library ieee;
use ieee.std_logic_1164.all;

package BOARD_ROM_VHDL_INIT is
type memory is array(0 to 32767) of std_logic_vector(7 downto 0);
constant init_vals : memory := (
-- note that the last addresses, i.e., those past your last 
--   non-zero data, can be replaced with the below line 
--   (without the leading dashes)
--   others => X"00"

x"00",	-- Hex Addr	0000	0
x"00",	-- Hex Addr	0001	1
x"00",	-- Hex Addr	0002	2
x"00",	-- Hex Addr	0003	3
x"00",	-- Hex Addr	0004	4
x"00",	-- Hex Addr	0005	5
x"00",	-- Hex Addr	0006	6
x"00",	-- Hex Addr	0007	7
x"00",	-- Hex Addr	0008	8
x"00",	-- Hex Addr	0009	9
x"00",	-- Hex Addr	000A	10
x"00",	-- Hex Addr	000B	11
x"00",	-- Hex Addr	000C	12
x"00",	-- Hex Addr	000D	13
x"00",	-- Hex Addr	000E	14
x"00",	-- Hex Addr	000F	15
x"00",	-- Hex Addr	0010	16
x"00",	-- Hex Addr	0011	17
x"00",	-- Hex Addr	0012	18
x"00",	-- Hex Addr	0013	19
x"00",	-- Hex Addr	0014	20
x"00",	-- Hex Addr	0015	21
x"00",	-- Hex Addr	0016	22
x"00",	-- Hex Addr	0017	23
x"00",	-- Hex Addr	0018	24
x"00",	-- Hex Addr	0019	25
x"00",	-- Hex Addr	001A	26
x"00",	-- Hex Addr	001B	27
x"00",	-- Hex Addr	001C	28
x"00",	-- Hex Addr	001D	29
x"00",	-- Hex Addr	001E	30
x"00",	-- Hex Addr	001F	31
x"00",	-- Hex Addr	0020	32
x"00",	-- Hex Addr	0021	33
x"00",	-- Hex Addr	0022	34
x"00",	-- Hex Addr	0023	35
x"00",	-- Hex Addr	0024	36
x"00",	-- Hex Addr	0025	37
x"00",	-- Hex Addr	0026	38
x"00",	-- Hex Addr	0027	39
x"00",	-- Hex Addr	0028	40
x"00",	-- Hex Addr	0029	41
x"00",	-- Hex Addr	002A	42
x"00",	-- Hex Addr	002B	43
x"00",	-- Hex Addr	002C	44
x"00",	-- Hex Addr	002D	45
x"00",	-- Hex Addr	002E	46
x"00",	-- Hex Addr	002F	47
x"00",	-- Hex Addr	0030	48
x"00",	-- Hex Addr	0031	49
x"00",	-- Hex Addr	0032	50
x"00",	-- Hex Addr	0033	51
x"00",	-- Hex Addr	0034	52
x"00",	-- Hex Addr	0035	53
x"00",	-- Hex Addr	0036	54
x"00",	-- Hex Addr	0037	55
x"00",	-- Hex Addr	0038	56
x"00",	-- Hex Addr	0039	57
x"00",	-- Hex Addr	003A	58
x"00",	-- Hex Addr	003B	59
x"00",	-- Hex Addr	003C	60
x"00",	-- Hex Addr	003D	61
x"00",	-- Hex Addr	003E	62
x"00",	-- Hex Addr	003F	63
x"00",	-- Hex Addr	0040	64
x"00",	-- Hex Addr	0041	65
x"00",	-- Hex Addr	0042	66
x"00",	-- Hex Addr	0043	67
x"00",	-- Hex Addr	0044	68
x"00",	-- Hex Addr	0045	69
x"00",	-- Hex Addr	0046	70
x"00",	-- Hex Addr	0047	71
x"00",	-- Hex Addr	0048	72
x"00",	-- Hex Addr	0049	73
x"00",	-- Hex Addr	004A	74
x"00",	-- Hex Addr	004B	75
x"00",	-- Hex Addr	004C	76
x"00",	-- Hex Addr	004D	77
x"00",	-- Hex Addr	004E	78
x"00",	-- Hex Addr	004F	79
x"00",	-- Hex Addr	0050	80
x"00",	-- Hex Addr	0051	81
x"00",	-- Hex Addr	0052	82
x"00",	-- Hex Addr	0053	83
x"00",	-- Hex Addr	0054	84
x"00",	-- Hex Addr	0055	85
x"00",	-- Hex Addr	0056	86
x"00",	-- Hex Addr	0057	87
x"00",	-- Hex Addr	0058	88
x"00",	-- Hex Addr	0059	89
x"00",	-- Hex Addr	005A	90
x"00",	-- Hex Addr	005B	91
x"00",	-- Hex Addr	005C	92
x"00",	-- Hex Addr	005D	93
x"00",	-- Hex Addr	005E	94
x"00",	-- Hex Addr	005F	95
x"00",	-- Hex Addr	0060	96
x"00",	-- Hex Addr	0061	97
x"00",	-- Hex Addr	0062	98
x"00",	-- Hex Addr	0063	99
x"00",	-- Hex Addr	0064	100
x"00",	-- Hex Addr	0065	101
x"00",	-- Hex Addr	0066	102
x"00",	-- Hex Addr	0067	103
x"00",	-- Hex Addr	0068	104
x"00",	-- Hex Addr	0069	105
x"00",	-- Hex Addr	006A	106
x"00",	-- Hex Addr	006B	107
x"00",	-- Hex Addr	006C	108
x"00",	-- Hex Addr	006D	109
x"00",	-- Hex Addr	006E	110
x"00",	-- Hex Addr	006F	111
x"00",	-- Hex Addr	0070	112
x"00",	-- Hex Addr	0071	113
x"00",	-- Hex Addr	0072	114
x"00",	-- Hex Addr	0073	115
x"00",	-- Hex Addr	0074	116
x"00",	-- Hex Addr	0075	117
x"00",	-- Hex Addr	0076	118
x"00",	-- Hex Addr	0077	119
x"00",	-- Hex Addr	0078	120
x"00",	-- Hex Addr	0079	121
x"00",	-- Hex Addr	007A	122
x"00",	-- Hex Addr	007B	123
x"00",	-- Hex Addr	007C	124
x"00",	-- Hex Addr	007D	125
x"00",	-- Hex Addr	007E	126
x"00",	-- Hex Addr	007F	127
x"00",	-- Hex Addr	0080	128
x"00",	-- Hex Addr	0081	129
x"00",	-- Hex Addr	0082	130
x"00",	-- Hex Addr	0083	131
x"00",	-- Hex Addr	0084	132
x"00",	-- Hex Addr	0085	133
x"00",	-- Hex Addr	0086	134
x"00",	-- Hex Addr	0087	135
x"00",	-- Hex Addr	0088	136
x"00",	-- Hex Addr	0089	137
x"00",	-- Hex Addr	008A	138
x"00",	-- Hex Addr	008B	139
x"00",	-- Hex Addr	008C	140
x"00",	-- Hex Addr	008D	141
x"00",	-- Hex Addr	008E	142
x"00",	-- Hex Addr	008F	143
x"00",	-- Hex Addr	0090	144
x"00",	-- Hex Addr	0091	145
x"00",	-- Hex Addr	0092	146
x"00",	-- Hex Addr	0093	147
x"00",	-- Hex Addr	0094	148
x"00",	-- Hex Addr	0095	149
x"00",	-- Hex Addr	0096	150
x"00",	-- Hex Addr	0097	151
x"00",	-- Hex Addr	0098	152
x"00",	-- Hex Addr	0099	153
x"00",	-- Hex Addr	009A	154
x"00",	-- Hex Addr	009B	155
x"00",	-- Hex Addr	009C	156
x"00",	-- Hex Addr	009D	157
x"00",	-- Hex Addr	009E	158
x"00",	-- Hex Addr	009F	159
x"00",	-- Hex Addr	00A0	160
x"00",	-- Hex Addr	00A1	161
x"00",	-- Hex Addr	00A2	162
x"00",	-- Hex Addr	00A3	163
x"00",	-- Hex Addr	00A4	164
x"00",	-- Hex Addr	00A5	165
x"00",	-- Hex Addr	00A6	166
x"00",	-- Hex Addr	00A7	167
x"00",	-- Hex Addr	00A8	168
x"00",	-- Hex Addr	00A9	169
x"00",	-- Hex Addr	00AA	170
x"00",	-- Hex Addr	00AB	171
x"00",	-- Hex Addr	00AC	172
x"00",	-- Hex Addr	00AD	173
x"00",	-- Hex Addr	00AE	174
x"00",	-- Hex Addr	00AF	175
x"00",	-- Hex Addr	00B0	176
x"00",	-- Hex Addr	00B1	177
x"00",	-- Hex Addr	00B2	178
x"00",	-- Hex Addr	00B3	179
x"00",	-- Hex Addr	00B4	180
x"00",	-- Hex Addr	00B5	181
x"00",	-- Hex Addr	00B6	182
x"00",	-- Hex Addr	00B7	183
x"00",	-- Hex Addr	00B8	184
x"00",	-- Hex Addr	00B9	185
x"00",	-- Hex Addr	00BA	186
x"00",	-- Hex Addr	00BB	187
x"00",	-- Hex Addr	00BC	188
x"00",	-- Hex Addr	00BD	189
x"00",	-- Hex Addr	00BE	190
x"00",	-- Hex Addr	00BF	191
x"00",	-- Hex Addr	00C0	192
x"00",	-- Hex Addr	00C1	193
x"00",	-- Hex Addr	00C2	194
x"00",	-- Hex Addr	00C3	195
x"00",	-- Hex Addr	00C4	196
x"00",	-- Hex Addr	00C5	197
x"00",	-- Hex Addr	00C6	198
x"00",	-- Hex Addr	00C7	199
x"00",	-- Hex Addr	00C8	200
x"00",	-- Hex Addr	00C9	201
x"00",	-- Hex Addr	00CA	202
x"00",	-- Hex Addr	00CB	203
x"00",	-- Hex Addr	00CC	204
x"00",	-- Hex Addr	00CD	205
x"00",	-- Hex Addr	00CE	206
x"00",	-- Hex Addr	00CF	207
x"00",	-- Hex Addr	00D0	208
x"00",	-- Hex Addr	00D1	209
x"00",	-- Hex Addr	00D2	210
x"00",	-- Hex Addr	00D3	211
x"00",	-- Hex Addr	00D4	212
x"00",	-- Hex Addr	00D5	213
x"00",	-- Hex Addr	00D6	214
x"00",	-- Hex Addr	00D7	215
x"00",	-- Hex Addr	00D8	216
x"00",	-- Hex Addr	00D9	217
x"00",	-- Hex Addr	00DA	218
x"00",	-- Hex Addr	00DB	219
x"00",	-- Hex Addr	00DC	220
x"00",	-- Hex Addr	00DD	221
x"00",	-- Hex Addr	00DE	222
x"00",	-- Hex Addr	00DF	223
x"00",	-- Hex Addr	00E0	224
x"00",	-- Hex Addr	00E1	225
x"00",	-- Hex Addr	00E2	226
x"00",	-- Hex Addr	00E3	227
x"00",	-- Hex Addr	00E4	228
x"00",	-- Hex Addr	00E5	229
x"00",	-- Hex Addr	00E6	230
x"00",	-- Hex Addr	00E7	231
x"00",	-- Hex Addr	00E8	232
x"00",	-- Hex Addr	00E9	233
x"00",	-- Hex Addr	00EA	234
x"00",	-- Hex Addr	00EB	235
x"00",	-- Hex Addr	00EC	236
x"00",	-- Hex Addr	00ED	237
x"00",	-- Hex Addr	00EE	238
x"00",	-- Hex Addr	00EF	239
x"00",	-- Hex Addr	00F0	240
x"00",	-- Hex Addr	00F1	241
x"00",	-- Hex Addr	00F2	242
x"00",	-- Hex Addr	00F3	243
x"00",	-- Hex Addr	00F4	244
x"00",	-- Hex Addr	00F5	245
x"00",	-- Hex Addr	00F6	246
x"00",	-- Hex Addr	00F7	247
x"00",	-- Hex Addr	00F8	248
x"00",	-- Hex Addr	00F9	249
x"00",	-- Hex Addr	00FA	250
x"00",	-- Hex Addr	00FB	251
x"00",	-- Hex Addr	00FC	252
x"00",	-- Hex Addr	00FD	253
x"00",	-- Hex Addr	00FE	254
x"00",	-- Hex Addr	00FF	255
x"00",	-- Hex Addr	0100	256
x"00",	-- Hex Addr	0101	257
x"00",	-- Hex Addr	0102	258
x"00",	-- Hex Addr	0103	259
x"00",	-- Hex Addr	0104	260
x"00",	-- Hex Addr	0105	261
x"00",	-- Hex Addr	0106	262
x"00",	-- Hex Addr	0107	263
x"00",	-- Hex Addr	0108	264
x"00",	-- Hex Addr	0109	265
x"00",	-- Hex Addr	010A	266
x"00",	-- Hex Addr	010B	267
x"00",	-- Hex Addr	010C	268
x"00",	-- Hex Addr	010D	269
x"00",	-- Hex Addr	010E	270
x"00",	-- Hex Addr	010F	271
x"00",	-- Hex Addr	0110	272
x"00",	-- Hex Addr	0111	273
x"00",	-- Hex Addr	0112	274
x"00",	-- Hex Addr	0113	275
x"00",	-- Hex Addr	0114	276
x"00",	-- Hex Addr	0115	277
x"00",	-- Hex Addr	0116	278
x"00",	-- Hex Addr	0117	279
x"00",	-- Hex Addr	0118	280
x"00",	-- Hex Addr	0119	281
x"00",	-- Hex Addr	011A	282
x"00",	-- Hex Addr	011B	283
x"00",	-- Hex Addr	011C	284
x"00",	-- Hex Addr	011D	285
x"00",	-- Hex Addr	011E	286
x"00",	-- Hex Addr	011F	287
x"00",	-- Hex Addr	0120	288
x"00",	-- Hex Addr	0121	289
x"00",	-- Hex Addr	0122	290
x"00",	-- Hex Addr	0123	291
x"00",	-- Hex Addr	0124	292
x"00",	-- Hex Addr	0125	293
x"00",	-- Hex Addr	0126	294
x"00",	-- Hex Addr	0127	295
x"00",	-- Hex Addr	0128	296
x"00",	-- Hex Addr	0129	297
x"00",	-- Hex Addr	012A	298
x"00",	-- Hex Addr	012B	299
x"00",	-- Hex Addr	012C	300
x"00",	-- Hex Addr	012D	301
x"00",	-- Hex Addr	012E	302
x"00",	-- Hex Addr	012F	303
x"00",	-- Hex Addr	0130	304
x"00",	-- Hex Addr	0131	305
x"00",	-- Hex Addr	0132	306
x"00",	-- Hex Addr	0133	307
x"00",	-- Hex Addr	0134	308
x"00",	-- Hex Addr	0135	309
x"00",	-- Hex Addr	0136	310
x"00",	-- Hex Addr	0137	311
x"00",	-- Hex Addr	0138	312
x"00",	-- Hex Addr	0139	313
x"00",	-- Hex Addr	013A	314
x"00",	-- Hex Addr	013B	315
x"00",	-- Hex Addr	013C	316
x"00",	-- Hex Addr	013D	317
x"00",	-- Hex Addr	013E	318
x"00",	-- Hex Addr	013F	319
x"00",	-- Hex Addr	0140	320
x"00",	-- Hex Addr	0141	321
x"00",	-- Hex Addr	0142	322
x"00",	-- Hex Addr	0143	323
x"00",	-- Hex Addr	0144	324
x"00",	-- Hex Addr	0145	325
x"00",	-- Hex Addr	0146	326
x"00",	-- Hex Addr	0147	327
x"00",	-- Hex Addr	0148	328
x"00",	-- Hex Addr	0149	329
x"00",	-- Hex Addr	014A	330
x"00",	-- Hex Addr	014B	331
x"00",	-- Hex Addr	014C	332
x"00",	-- Hex Addr	014D	333
x"00",	-- Hex Addr	014E	334
x"00",	-- Hex Addr	014F	335
x"00",	-- Hex Addr	0150	336
x"00",	-- Hex Addr	0151	337
x"00",	-- Hex Addr	0152	338
x"00",	-- Hex Addr	0153	339
x"00",	-- Hex Addr	0154	340
x"00",	-- Hex Addr	0155	341
x"00",	-- Hex Addr	0156	342
x"00",	-- Hex Addr	0157	343
x"00",	-- Hex Addr	0158	344
x"00",	-- Hex Addr	0159	345
x"00",	-- Hex Addr	015A	346
x"00",	-- Hex Addr	015B	347
x"00",	-- Hex Addr	015C	348
x"00",	-- Hex Addr	015D	349
x"00",	-- Hex Addr	015E	350
x"00",	-- Hex Addr	015F	351
x"00",	-- Hex Addr	0160	352
x"00",	-- Hex Addr	0161	353
x"00",	-- Hex Addr	0162	354
x"00",	-- Hex Addr	0163	355
x"00",	-- Hex Addr	0164	356
x"00",	-- Hex Addr	0165	357
x"00",	-- Hex Addr	0166	358
x"00",	-- Hex Addr	0167	359
x"00",	-- Hex Addr	0168	360
x"00",	-- Hex Addr	0169	361
x"00",	-- Hex Addr	016A	362
x"00",	-- Hex Addr	016B	363
x"00",	-- Hex Addr	016C	364
x"00",	-- Hex Addr	016D	365
x"00",	-- Hex Addr	016E	366
x"00",	-- Hex Addr	016F	367
x"00",	-- Hex Addr	0170	368
x"00",	-- Hex Addr	0171	369
x"00",	-- Hex Addr	0172	370
x"00",	-- Hex Addr	0173	371
x"00",	-- Hex Addr	0174	372
x"00",	-- Hex Addr	0175	373
x"00",	-- Hex Addr	0176	374
x"00",	-- Hex Addr	0177	375
x"00",	-- Hex Addr	0178	376
x"00",	-- Hex Addr	0179	377
x"00",	-- Hex Addr	017A	378
x"00",	-- Hex Addr	017B	379
x"00",	-- Hex Addr	017C	380
x"00",	-- Hex Addr	017D	381
x"00",	-- Hex Addr	017E	382
x"00",	-- Hex Addr	017F	383
x"00",	-- Hex Addr	0180	384
x"00",	-- Hex Addr	0181	385
x"00",	-- Hex Addr	0182	386
x"00",	-- Hex Addr	0183	387
x"00",	-- Hex Addr	0184	388
x"00",	-- Hex Addr	0185	389
x"00",	-- Hex Addr	0186	390
x"00",	-- Hex Addr	0187	391
x"00",	-- Hex Addr	0188	392
x"00",	-- Hex Addr	0189	393
x"00",	-- Hex Addr	018A	394
x"00",	-- Hex Addr	018B	395
x"00",	-- Hex Addr	018C	396
x"00",	-- Hex Addr	018D	397
x"00",	-- Hex Addr	018E	398
x"00",	-- Hex Addr	018F	399
x"00",	-- Hex Addr	0190	400
x"00",	-- Hex Addr	0191	401
x"00",	-- Hex Addr	0192	402
x"00",	-- Hex Addr	0193	403
x"00",	-- Hex Addr	0194	404
x"00",	-- Hex Addr	0195	405
x"00",	-- Hex Addr	0196	406
x"00",	-- Hex Addr	0197	407
x"00",	-- Hex Addr	0198	408
x"00",	-- Hex Addr	0199	409
x"00",	-- Hex Addr	019A	410
x"00",	-- Hex Addr	019B	411
x"00",	-- Hex Addr	019C	412
x"00",	-- Hex Addr	019D	413
x"00",	-- Hex Addr	019E	414
x"00",	-- Hex Addr	019F	415
x"00",	-- Hex Addr	01A0	416
x"00",	-- Hex Addr	01A1	417
x"00",	-- Hex Addr	01A2	418
x"00",	-- Hex Addr	01A3	419
x"00",	-- Hex Addr	01A4	420
x"00",	-- Hex Addr	01A5	421
x"00",	-- Hex Addr	01A6	422
x"00",	-- Hex Addr	01A7	423
x"00",	-- Hex Addr	01A8	424
x"00",	-- Hex Addr	01A9	425
x"00",	-- Hex Addr	01AA	426
x"00",	-- Hex Addr	01AB	427
x"00",	-- Hex Addr	01AC	428
x"00",	-- Hex Addr	01AD	429
x"00",	-- Hex Addr	01AE	430
x"00",	-- Hex Addr	01AF	431
x"00",	-- Hex Addr	01B0	432
x"00",	-- Hex Addr	01B1	433
x"00",	-- Hex Addr	01B2	434
x"00",	-- Hex Addr	01B3	435
x"00",	-- Hex Addr	01B4	436
x"00",	-- Hex Addr	01B5	437
x"00",	-- Hex Addr	01B6	438
x"00",	-- Hex Addr	01B7	439
x"00",	-- Hex Addr	01B8	440
x"00",	-- Hex Addr	01B9	441
x"00",	-- Hex Addr	01BA	442
x"00",	-- Hex Addr	01BB	443
x"00",	-- Hex Addr	01BC	444
x"00",	-- Hex Addr	01BD	445
x"00",	-- Hex Addr	01BE	446
x"00",	-- Hex Addr	01BF	447
x"00",	-- Hex Addr	01C0	448
x"00",	-- Hex Addr	01C1	449
x"00",	-- Hex Addr	01C2	450
x"00",	-- Hex Addr	01C3	451
x"00",	-- Hex Addr	01C4	452
x"00",	-- Hex Addr	01C5	453
x"00",	-- Hex Addr	01C6	454
x"00",	-- Hex Addr	01C7	455
x"00",	-- Hex Addr	01C8	456
x"00",	-- Hex Addr	01C9	457
x"00",	-- Hex Addr	01CA	458
x"00",	-- Hex Addr	01CB	459
x"00",	-- Hex Addr	01CC	460
x"00",	-- Hex Addr	01CD	461
x"00",	-- Hex Addr	01CE	462
x"00",	-- Hex Addr	01CF	463
x"00",	-- Hex Addr	01D0	464
x"00",	-- Hex Addr	01D1	465
x"00",	-- Hex Addr	01D2	466
x"00",	-- Hex Addr	01D3	467
x"00",	-- Hex Addr	01D4	468
x"00",	-- Hex Addr	01D5	469
x"00",	-- Hex Addr	01D6	470
x"00",	-- Hex Addr	01D7	471
x"00",	-- Hex Addr	01D8	472
x"00",	-- Hex Addr	01D9	473
x"00",	-- Hex Addr	01DA	474
x"00",	-- Hex Addr	01DB	475
x"00",	-- Hex Addr	01DC	476
x"00",	-- Hex Addr	01DD	477
x"00",	-- Hex Addr	01DE	478
x"00",	-- Hex Addr	01DF	479
x"00",	-- Hex Addr	01E0	480
x"00",	-- Hex Addr	01E1	481
x"00",	-- Hex Addr	01E2	482
x"00",	-- Hex Addr	01E3	483
x"00",	-- Hex Addr	01E4	484
x"00",	-- Hex Addr	01E5	485
x"00",	-- Hex Addr	01E6	486
x"00",	-- Hex Addr	01E7	487
x"00",	-- Hex Addr	01E8	488
x"00",	-- Hex Addr	01E9	489
x"00",	-- Hex Addr	01EA	490
x"00",	-- Hex Addr	01EB	491
x"00",	-- Hex Addr	01EC	492
x"00",	-- Hex Addr	01ED	493
x"00",	-- Hex Addr	01EE	494
x"00",	-- Hex Addr	01EF	495
x"00",	-- Hex Addr	01F0	496
x"00",	-- Hex Addr	01F1	497
x"00",	-- Hex Addr	01F2	498
x"00",	-- Hex Addr	01F3	499
x"00",	-- Hex Addr	01F4	500
x"00",	-- Hex Addr	01F5	501
x"00",	-- Hex Addr	01F6	502
x"00",	-- Hex Addr	01F7	503
x"00",	-- Hex Addr	01F8	504
x"00",	-- Hex Addr	01F9	505
x"00",	-- Hex Addr	01FA	506
x"00",	-- Hex Addr	01FB	507
x"00",	-- Hex Addr	01FC	508
x"00",	-- Hex Addr	01FD	509
x"00",	-- Hex Addr	01FE	510
x"00",	-- Hex Addr	01FF	511
x"00",	-- Hex Addr	0200	512
x"00",	-- Hex Addr	0201	513
x"00",	-- Hex Addr	0202	514
x"00",	-- Hex Addr	0203	515
x"00",	-- Hex Addr	0204	516
x"00",	-- Hex Addr	0205	517
x"00",	-- Hex Addr	0206	518
x"00",	-- Hex Addr	0207	519
x"00",	-- Hex Addr	0208	520
x"00",	-- Hex Addr	0209	521
x"00",	-- Hex Addr	020A	522
x"00",	-- Hex Addr	020B	523
x"00",	-- Hex Addr	020C	524
x"00",	-- Hex Addr	020D	525
x"00",	-- Hex Addr	020E	526
x"00",	-- Hex Addr	020F	527
x"00",	-- Hex Addr	0210	528
x"00",	-- Hex Addr	0211	529
x"00",	-- Hex Addr	0212	530
x"00",	-- Hex Addr	0213	531
x"00",	-- Hex Addr	0214	532
x"00",	-- Hex Addr	0215	533
x"00",	-- Hex Addr	0216	534
x"00",	-- Hex Addr	0217	535
x"00",	-- Hex Addr	0218	536
x"00",	-- Hex Addr	0219	537
x"00",	-- Hex Addr	021A	538
x"00",	-- Hex Addr	021B	539
x"00",	-- Hex Addr	021C	540
x"00",	-- Hex Addr	021D	541
x"00",	-- Hex Addr	021E	542
x"00",	-- Hex Addr	021F	543
x"00",	-- Hex Addr	0220	544
x"00",	-- Hex Addr	0221	545
x"00",	-- Hex Addr	0222	546
x"00",	-- Hex Addr	0223	547
x"00",	-- Hex Addr	0224	548
x"00",	-- Hex Addr	0225	549
x"00",	-- Hex Addr	0226	550
x"00",	-- Hex Addr	0227	551
x"00",	-- Hex Addr	0228	552
x"00",	-- Hex Addr	0229	553
x"00",	-- Hex Addr	022A	554
x"00",	-- Hex Addr	022B	555
x"00",	-- Hex Addr	022C	556
x"00",	-- Hex Addr	022D	557
x"00",	-- Hex Addr	022E	558
x"00",	-- Hex Addr	022F	559
x"00",	-- Hex Addr	0230	560
x"00",	-- Hex Addr	0231	561
x"00",	-- Hex Addr	0232	562
x"00",	-- Hex Addr	0233	563
x"00",	-- Hex Addr	0234	564
x"00",	-- Hex Addr	0235	565
x"00",	-- Hex Addr	0236	566
x"00",	-- Hex Addr	0237	567
x"00",	-- Hex Addr	0238	568
x"00",	-- Hex Addr	0239	569
x"00",	-- Hex Addr	023A	570
x"00",	-- Hex Addr	023B	571
x"00",	-- Hex Addr	023C	572
x"00",	-- Hex Addr	023D	573
x"00",	-- Hex Addr	023E	574
x"00",	-- Hex Addr	023F	575
x"00",	-- Hex Addr	0240	576
x"00",	-- Hex Addr	0241	577
x"00",	-- Hex Addr	0242	578
x"00",	-- Hex Addr	0243	579
x"00",	-- Hex Addr	0244	580
x"00",	-- Hex Addr	0245	581
x"00",	-- Hex Addr	0246	582
x"00",	-- Hex Addr	0247	583
x"00",	-- Hex Addr	0248	584
x"00",	-- Hex Addr	0249	585
x"00",	-- Hex Addr	024A	586
x"00",	-- Hex Addr	024B	587
x"00",	-- Hex Addr	024C	588
x"00",	-- Hex Addr	024D	589
x"00",	-- Hex Addr	024E	590
x"00",	-- Hex Addr	024F	591
x"00",	-- Hex Addr	0250	592
x"00",	-- Hex Addr	0251	593
x"00",	-- Hex Addr	0252	594
x"00",	-- Hex Addr	0253	595
x"00",	-- Hex Addr	0254	596
x"00",	-- Hex Addr	0255	597
x"00",	-- Hex Addr	0256	598
x"00",	-- Hex Addr	0257	599
x"00",	-- Hex Addr	0258	600
x"00",	-- Hex Addr	0259	601
x"00",	-- Hex Addr	025A	602
x"00",	-- Hex Addr	025B	603
x"00",	-- Hex Addr	025C	604
x"00",	-- Hex Addr	025D	605
x"00",	-- Hex Addr	025E	606
x"00",	-- Hex Addr	025F	607
x"00",	-- Hex Addr	0260	608
x"00",	-- Hex Addr	0261	609
x"00",	-- Hex Addr	0262	610
x"00",	-- Hex Addr	0263	611
x"00",	-- Hex Addr	0264	612
x"00",	-- Hex Addr	0265	613
x"00",	-- Hex Addr	0266	614
x"00",	-- Hex Addr	0267	615
x"00",	-- Hex Addr	0268	616
x"00",	-- Hex Addr	0269	617
x"00",	-- Hex Addr	026A	618
x"00",	-- Hex Addr	026B	619
x"00",	-- Hex Addr	026C	620
x"00",	-- Hex Addr	026D	621
x"00",	-- Hex Addr	026E	622
x"00",	-- Hex Addr	026F	623
x"00",	-- Hex Addr	0270	624
x"00",	-- Hex Addr	0271	625
x"00",	-- Hex Addr	0272	626
x"00",	-- Hex Addr	0273	627
x"00",	-- Hex Addr	0274	628
x"00",	-- Hex Addr	0275	629
x"00",	-- Hex Addr	0276	630
x"00",	-- Hex Addr	0277	631
x"00",	-- Hex Addr	0278	632
x"00",	-- Hex Addr	0279	633
x"00",	-- Hex Addr	027A	634
x"00",	-- Hex Addr	027B	635
x"00",	-- Hex Addr	027C	636
x"00",	-- Hex Addr	027D	637
x"00",	-- Hex Addr	027E	638
x"00",	-- Hex Addr	027F	639
x"00",	-- Hex Addr	0280	640
x"00",	-- Hex Addr	0281	641
x"00",	-- Hex Addr	0282	642
x"00",	-- Hex Addr	0283	643
x"00",	-- Hex Addr	0284	644
x"00",	-- Hex Addr	0285	645
x"00",	-- Hex Addr	0286	646
x"00",	-- Hex Addr	0287	647
x"00",	-- Hex Addr	0288	648
x"00",	-- Hex Addr	0289	649
x"00",	-- Hex Addr	028A	650
x"00",	-- Hex Addr	028B	651
x"00",	-- Hex Addr	028C	652
x"00",	-- Hex Addr	028D	653
x"00",	-- Hex Addr	028E	654
x"00",	-- Hex Addr	028F	655
x"00",	-- Hex Addr	0290	656
x"00",	-- Hex Addr	0291	657
x"00",	-- Hex Addr	0292	658
x"00",	-- Hex Addr	0293	659
x"00",	-- Hex Addr	0294	660
x"00",	-- Hex Addr	0295	661
x"00",	-- Hex Addr	0296	662
x"00",	-- Hex Addr	0297	663
x"00",	-- Hex Addr	0298	664
x"00",	-- Hex Addr	0299	665
x"00",	-- Hex Addr	029A	666
x"00",	-- Hex Addr	029B	667
x"00",	-- Hex Addr	029C	668
x"00",	-- Hex Addr	029D	669
x"00",	-- Hex Addr	029E	670
x"00",	-- Hex Addr	029F	671
x"00",	-- Hex Addr	02A0	672
x"00",	-- Hex Addr	02A1	673
x"00",	-- Hex Addr	02A2	674
x"00",	-- Hex Addr	02A3	675
x"00",	-- Hex Addr	02A4	676
x"00",	-- Hex Addr	02A5	677
x"00",	-- Hex Addr	02A6	678
x"00",	-- Hex Addr	02A7	679
x"00",	-- Hex Addr	02A8	680
x"00",	-- Hex Addr	02A9	681
x"00",	-- Hex Addr	02AA	682
x"00",	-- Hex Addr	02AB	683
x"00",	-- Hex Addr	02AC	684
x"00",	-- Hex Addr	02AD	685
x"00",	-- Hex Addr	02AE	686
x"00",	-- Hex Addr	02AF	687
x"00",	-- Hex Addr	02B0	688
x"00",	-- Hex Addr	02B1	689
x"00",	-- Hex Addr	02B2	690
x"00",	-- Hex Addr	02B3	691
x"00",	-- Hex Addr	02B4	692
x"00",	-- Hex Addr	02B5	693
x"00",	-- Hex Addr	02B6	694
x"00",	-- Hex Addr	02B7	695
x"00",	-- Hex Addr	02B8	696
x"00",	-- Hex Addr	02B9	697
x"00",	-- Hex Addr	02BA	698
x"00",	-- Hex Addr	02BB	699
x"00",	-- Hex Addr	02BC	700
x"00",	-- Hex Addr	02BD	701
x"00",	-- Hex Addr	02BE	702
x"00",	-- Hex Addr	02BF	703
x"00",	-- Hex Addr	02C0	704
x"00",	-- Hex Addr	02C1	705
x"00",	-- Hex Addr	02C2	706
x"00",	-- Hex Addr	02C3	707
x"00",	-- Hex Addr	02C4	708
x"00",	-- Hex Addr	02C5	709
x"00",	-- Hex Addr	02C6	710
x"00",	-- Hex Addr	02C7	711
x"00",	-- Hex Addr	02C8	712
x"00",	-- Hex Addr	02C9	713
x"00",	-- Hex Addr	02CA	714
x"00",	-- Hex Addr	02CB	715
x"00",	-- Hex Addr	02CC	716
x"00",	-- Hex Addr	02CD	717
x"00",	-- Hex Addr	02CE	718
x"00",	-- Hex Addr	02CF	719
x"00",	-- Hex Addr	02D0	720
x"00",	-- Hex Addr	02D1	721
x"00",	-- Hex Addr	02D2	722
x"00",	-- Hex Addr	02D3	723
x"00",	-- Hex Addr	02D4	724
x"00",	-- Hex Addr	02D5	725
x"00",	-- Hex Addr	02D6	726
x"00",	-- Hex Addr	02D7	727
x"00",	-- Hex Addr	02D8	728
x"00",	-- Hex Addr	02D9	729
x"00",	-- Hex Addr	02DA	730
x"00",	-- Hex Addr	02DB	731
x"00",	-- Hex Addr	02DC	732
x"00",	-- Hex Addr	02DD	733
x"00",	-- Hex Addr	02DE	734
x"00",	-- Hex Addr	02DF	735
x"00",	-- Hex Addr	02E0	736
x"00",	-- Hex Addr	02E1	737
x"00",	-- Hex Addr	02E2	738
x"00",	-- Hex Addr	02E3	739
x"00",	-- Hex Addr	02E4	740
x"00",	-- Hex Addr	02E5	741
x"00",	-- Hex Addr	02E6	742
x"00",	-- Hex Addr	02E7	743
x"00",	-- Hex Addr	02E8	744
x"00",	-- Hex Addr	02E9	745
x"00",	-- Hex Addr	02EA	746
x"00",	-- Hex Addr	02EB	747
x"00",	-- Hex Addr	02EC	748
x"00",	-- Hex Addr	02ED	749
x"00",	-- Hex Addr	02EE	750
x"00",	-- Hex Addr	02EF	751
x"00",	-- Hex Addr	02F0	752
x"00",	-- Hex Addr	02F1	753
x"00",	-- Hex Addr	02F2	754
x"00",	-- Hex Addr	02F3	755
x"00",	-- Hex Addr	02F4	756
x"00",	-- Hex Addr	02F5	757
x"00",	-- Hex Addr	02F6	758
x"00",	-- Hex Addr	02F7	759
x"00",	-- Hex Addr	02F8	760
x"00",	-- Hex Addr	02F9	761
x"00",	-- Hex Addr	02FA	762
x"00",	-- Hex Addr	02FB	763
x"00",	-- Hex Addr	02FC	764
x"00",	-- Hex Addr	02FD	765
x"00",	-- Hex Addr	02FE	766
x"00",	-- Hex Addr	02FF	767
x"00",	-- Hex Addr	0300	768
x"00",	-- Hex Addr	0301	769
x"00",	-- Hex Addr	0302	770
x"00",	-- Hex Addr	0303	771
x"00",	-- Hex Addr	0304	772
x"00",	-- Hex Addr	0305	773
x"00",	-- Hex Addr	0306	774
x"00",	-- Hex Addr	0307	775
x"00",	-- Hex Addr	0308	776
x"00",	-- Hex Addr	0309	777
x"00",	-- Hex Addr	030A	778
x"00",	-- Hex Addr	030B	779
x"00",	-- Hex Addr	030C	780
x"00",	-- Hex Addr	030D	781
x"00",	-- Hex Addr	030E	782
x"00",	-- Hex Addr	030F	783
x"00",	-- Hex Addr	0310	784
x"00",	-- Hex Addr	0311	785
x"00",	-- Hex Addr	0312	786
x"00",	-- Hex Addr	0313	787
x"00",	-- Hex Addr	0314	788
x"00",	-- Hex Addr	0315	789
x"00",	-- Hex Addr	0316	790
x"00",	-- Hex Addr	0317	791
x"00",	-- Hex Addr	0318	792
x"00",	-- Hex Addr	0319	793
x"00",	-- Hex Addr	031A	794
x"00",	-- Hex Addr	031B	795
x"00",	-- Hex Addr	031C	796
x"00",	-- Hex Addr	031D	797
x"00",	-- Hex Addr	031E	798
x"00",	-- Hex Addr	031F	799
x"00",	-- Hex Addr	0320	800
x"00",	-- Hex Addr	0321	801
x"00",	-- Hex Addr	0322	802
x"00",	-- Hex Addr	0323	803
x"00",	-- Hex Addr	0324	804
x"00",	-- Hex Addr	0325	805
x"00",	-- Hex Addr	0326	806
x"00",	-- Hex Addr	0327	807
x"00",	-- Hex Addr	0328	808
x"00",	-- Hex Addr	0329	809
x"00",	-- Hex Addr	032A	810
x"00",	-- Hex Addr	032B	811
x"00",	-- Hex Addr	032C	812
x"00",	-- Hex Addr	032D	813
x"00",	-- Hex Addr	032E	814
x"00",	-- Hex Addr	032F	815
x"00",	-- Hex Addr	0330	816
x"00",	-- Hex Addr	0331	817
x"00",	-- Hex Addr	0332	818
x"00",	-- Hex Addr	0333	819
x"00",	-- Hex Addr	0334	820
x"00",	-- Hex Addr	0335	821
x"00",	-- Hex Addr	0336	822
x"00",	-- Hex Addr	0337	823
x"00",	-- Hex Addr	0338	824
x"00",	-- Hex Addr	0339	825
x"00",	-- Hex Addr	033A	826
x"00",	-- Hex Addr	033B	827
x"00",	-- Hex Addr	033C	828
x"00",	-- Hex Addr	033D	829
x"00",	-- Hex Addr	033E	830
x"00",	-- Hex Addr	033F	831
x"00",	-- Hex Addr	0340	832
x"00",	-- Hex Addr	0341	833
x"00",	-- Hex Addr	0342	834
x"00",	-- Hex Addr	0343	835
x"00",	-- Hex Addr	0344	836
x"00",	-- Hex Addr	0345	837
x"00",	-- Hex Addr	0346	838
x"00",	-- Hex Addr	0347	839
x"00",	-- Hex Addr	0348	840
x"00",	-- Hex Addr	0349	841
x"00",	-- Hex Addr	034A	842
x"00",	-- Hex Addr	034B	843
x"00",	-- Hex Addr	034C	844
x"00",	-- Hex Addr	034D	845
x"00",	-- Hex Addr	034E	846
x"00",	-- Hex Addr	034F	847
x"00",	-- Hex Addr	0350	848
x"00",	-- Hex Addr	0351	849
x"00",	-- Hex Addr	0352	850
x"00",	-- Hex Addr	0353	851
x"00",	-- Hex Addr	0354	852
x"00",	-- Hex Addr	0355	853
x"00",	-- Hex Addr	0356	854
x"00",	-- Hex Addr	0357	855
x"00",	-- Hex Addr	0358	856
x"00",	-- Hex Addr	0359	857
x"00",	-- Hex Addr	035A	858
x"00",	-- Hex Addr	035B	859
x"00",	-- Hex Addr	035C	860
x"00",	-- Hex Addr	035D	861
x"00",	-- Hex Addr	035E	862
x"00",	-- Hex Addr	035F	863
x"00",	-- Hex Addr	0360	864
x"00",	-- Hex Addr	0361	865
x"00",	-- Hex Addr	0362	866
x"00",	-- Hex Addr	0363	867
x"00",	-- Hex Addr	0364	868
x"00",	-- Hex Addr	0365	869
x"00",	-- Hex Addr	0366	870
x"00",	-- Hex Addr	0367	871
x"00",	-- Hex Addr	0368	872
x"00",	-- Hex Addr	0369	873
x"00",	-- Hex Addr	036A	874
x"00",	-- Hex Addr	036B	875
x"00",	-- Hex Addr	036C	876
x"00",	-- Hex Addr	036D	877
x"00",	-- Hex Addr	036E	878
x"00",	-- Hex Addr	036F	879
x"00",	-- Hex Addr	0370	880
x"00",	-- Hex Addr	0371	881
x"00",	-- Hex Addr	0372	882
x"00",	-- Hex Addr	0373	883
x"00",	-- Hex Addr	0374	884
x"00",	-- Hex Addr	0375	885
x"00",	-- Hex Addr	0376	886
x"00",	-- Hex Addr	0377	887
x"00",	-- Hex Addr	0378	888
x"00",	-- Hex Addr	0379	889
x"00",	-- Hex Addr	037A	890
x"00",	-- Hex Addr	037B	891
x"00",	-- Hex Addr	037C	892
x"00",	-- Hex Addr	037D	893
x"00",	-- Hex Addr	037E	894
x"00",	-- Hex Addr	037F	895
x"00",	-- Hex Addr	0380	896
x"00",	-- Hex Addr	0381	897
x"00",	-- Hex Addr	0382	898
x"00",	-- Hex Addr	0383	899
x"00",	-- Hex Addr	0384	900
x"00",	-- Hex Addr	0385	901
x"00",	-- Hex Addr	0386	902
x"00",	-- Hex Addr	0387	903
x"00",	-- Hex Addr	0388	904
x"00",	-- Hex Addr	0389	905
x"00",	-- Hex Addr	038A	906
x"00",	-- Hex Addr	038B	907
x"00",	-- Hex Addr	038C	908
x"00",	-- Hex Addr	038D	909
x"00",	-- Hex Addr	038E	910
x"00",	-- Hex Addr	038F	911
x"00",	-- Hex Addr	0390	912
x"00",	-- Hex Addr	0391	913
x"00",	-- Hex Addr	0392	914
x"00",	-- Hex Addr	0393	915
x"00",	-- Hex Addr	0394	916
x"00",	-- Hex Addr	0395	917
x"00",	-- Hex Addr	0396	918
x"00",	-- Hex Addr	0397	919
x"00",	-- Hex Addr	0398	920
x"00",	-- Hex Addr	0399	921
x"00",	-- Hex Addr	039A	922
x"00",	-- Hex Addr	039B	923
x"00",	-- Hex Addr	039C	924
x"00",	-- Hex Addr	039D	925
x"00",	-- Hex Addr	039E	926
x"00",	-- Hex Addr	039F	927
x"00",	-- Hex Addr	03A0	928
x"00",	-- Hex Addr	03A1	929
x"00",	-- Hex Addr	03A2	930
x"00",	-- Hex Addr	03A3	931
x"00",	-- Hex Addr	03A4	932
x"00",	-- Hex Addr	03A5	933
x"00",	-- Hex Addr	03A6	934
x"00",	-- Hex Addr	03A7	935
x"00",	-- Hex Addr	03A8	936
x"00",	-- Hex Addr	03A9	937
x"00",	-- Hex Addr	03AA	938
x"00",	-- Hex Addr	03AB	939
x"00",	-- Hex Addr	03AC	940
x"00",	-- Hex Addr	03AD	941
x"00",	-- Hex Addr	03AE	942
x"00",	-- Hex Addr	03AF	943
x"00",	-- Hex Addr	03B0	944
x"00",	-- Hex Addr	03B1	945
x"00",	-- Hex Addr	03B2	946
x"00",	-- Hex Addr	03B3	947
x"00",	-- Hex Addr	03B4	948
x"00",	-- Hex Addr	03B5	949
x"00",	-- Hex Addr	03B6	950
x"00",	-- Hex Addr	03B7	951
x"00",	-- Hex Addr	03B8	952
x"00",	-- Hex Addr	03B9	953
x"00",	-- Hex Addr	03BA	954
x"00",	-- Hex Addr	03BB	955
x"00",	-- Hex Addr	03BC	956
x"00",	-- Hex Addr	03BD	957
x"00",	-- Hex Addr	03BE	958
x"00",	-- Hex Addr	03BF	959
x"00",	-- Hex Addr	03C0	960
x"00",	-- Hex Addr	03C1	961
x"00",	-- Hex Addr	03C2	962
x"00",	-- Hex Addr	03C3	963
x"00",	-- Hex Addr	03C4	964
x"00",	-- Hex Addr	03C5	965
x"00",	-- Hex Addr	03C6	966
x"00",	-- Hex Addr	03C7	967
x"00",	-- Hex Addr	03C8	968
x"00",	-- Hex Addr	03C9	969
x"00",	-- Hex Addr	03CA	970
x"00",	-- Hex Addr	03CB	971
x"00",	-- Hex Addr	03CC	972
x"00",	-- Hex Addr	03CD	973
x"00",	-- Hex Addr	03CE	974
x"00",	-- Hex Addr	03CF	975
x"00",	-- Hex Addr	03D0	976
x"00",	-- Hex Addr	03D1	977
x"00",	-- Hex Addr	03D2	978
x"00",	-- Hex Addr	03D3	979
x"00",	-- Hex Addr	03D4	980
x"00",	-- Hex Addr	03D5	981
x"00",	-- Hex Addr	03D6	982
x"00",	-- Hex Addr	03D7	983
x"00",	-- Hex Addr	03D8	984
x"00",	-- Hex Addr	03D9	985
x"00",	-- Hex Addr	03DA	986
x"00",	-- Hex Addr	03DB	987
x"00",	-- Hex Addr	03DC	988
x"00",	-- Hex Addr	03DD	989
x"00",	-- Hex Addr	03DE	990
x"00",	-- Hex Addr	03DF	991
x"00",	-- Hex Addr	03E0	992
x"00",	-- Hex Addr	03E1	993
x"00",	-- Hex Addr	03E2	994
x"00",	-- Hex Addr	03E3	995
x"00",	-- Hex Addr	03E4	996
x"00",	-- Hex Addr	03E5	997
x"00",	-- Hex Addr	03E6	998
x"00",	-- Hex Addr	03E7	999
x"00",	-- Hex Addr	03E8	1000
x"00",	-- Hex Addr	03E9	1001
x"00",	-- Hex Addr	03EA	1002
x"00",	-- Hex Addr	03EB	1003
x"00",	-- Hex Addr	03EC	1004
x"00",	-- Hex Addr	03ED	1005
x"00",	-- Hex Addr	03EE	1006
x"00",	-- Hex Addr	03EF	1007
x"00",	-- Hex Addr	03F0	1008
x"00",	-- Hex Addr	03F1	1009
x"00",	-- Hex Addr	03F2	1010
x"00",	-- Hex Addr	03F3	1011
x"00",	-- Hex Addr	03F4	1012
x"00",	-- Hex Addr	03F5	1013
x"00",	-- Hex Addr	03F6	1014
x"00",	-- Hex Addr	03F7	1015
x"00",	-- Hex Addr	03F8	1016
x"00",	-- Hex Addr	03F9	1017
x"00",	-- Hex Addr	03FA	1018
x"00",	-- Hex Addr	03FB	1019
x"00",	-- Hex Addr	03FC	1020
x"00",	-- Hex Addr	03FD	1021
x"00",	-- Hex Addr	03FE	1022
x"00",	-- Hex Addr	03FF	1023
x"00",	-- Hex Addr	0400	1024
x"00",	-- Hex Addr	0401	1025
x"00",	-- Hex Addr	0402	1026
x"00",	-- Hex Addr	0403	1027
x"00",	-- Hex Addr	0404	1028
x"00",	-- Hex Addr	0405	1029
x"00",	-- Hex Addr	0406	1030
x"00",	-- Hex Addr	0407	1031
x"00",	-- Hex Addr	0408	1032
x"00",	-- Hex Addr	0409	1033
x"00",	-- Hex Addr	040A	1034
x"00",	-- Hex Addr	040B	1035
x"00",	-- Hex Addr	040C	1036
x"00",	-- Hex Addr	040D	1037
x"00",	-- Hex Addr	040E	1038
x"00",	-- Hex Addr	040F	1039
x"00",	-- Hex Addr	0410	1040
x"00",	-- Hex Addr	0411	1041
x"00",	-- Hex Addr	0412	1042
x"00",	-- Hex Addr	0413	1043
x"00",	-- Hex Addr	0414	1044
x"00",	-- Hex Addr	0415	1045
x"00",	-- Hex Addr	0416	1046
x"00",	-- Hex Addr	0417	1047
x"00",	-- Hex Addr	0418	1048
x"00",	-- Hex Addr	0419	1049
x"00",	-- Hex Addr	041A	1050
x"00",	-- Hex Addr	041B	1051
x"00",	-- Hex Addr	041C	1052
x"00",	-- Hex Addr	041D	1053
x"00",	-- Hex Addr	041E	1054
x"00",	-- Hex Addr	041F	1055
x"00",	-- Hex Addr	0420	1056
x"00",	-- Hex Addr	0421	1057
x"00",	-- Hex Addr	0422	1058
x"00",	-- Hex Addr	0423	1059
x"00",	-- Hex Addr	0424	1060
x"00",	-- Hex Addr	0425	1061
x"00",	-- Hex Addr	0426	1062
x"00",	-- Hex Addr	0427	1063
x"00",	-- Hex Addr	0428	1064
x"00",	-- Hex Addr	0429	1065
x"00",	-- Hex Addr	042A	1066
x"00",	-- Hex Addr	042B	1067
x"00",	-- Hex Addr	042C	1068
x"00",	-- Hex Addr	042D	1069
x"00",	-- Hex Addr	042E	1070
x"00",	-- Hex Addr	042F	1071
x"00",	-- Hex Addr	0430	1072
x"00",	-- Hex Addr	0431	1073
x"00",	-- Hex Addr	0432	1074
x"00",	-- Hex Addr	0433	1075
x"00",	-- Hex Addr	0434	1076
x"00",	-- Hex Addr	0435	1077
x"00",	-- Hex Addr	0436	1078
x"00",	-- Hex Addr	0437	1079
x"00",	-- Hex Addr	0438	1080
x"00",	-- Hex Addr	0439	1081
x"00",	-- Hex Addr	043A	1082
x"00",	-- Hex Addr	043B	1083
x"00",	-- Hex Addr	043C	1084
x"00",	-- Hex Addr	043D	1085
x"00",	-- Hex Addr	043E	1086
x"00",	-- Hex Addr	043F	1087
x"00",	-- Hex Addr	0440	1088
x"00",	-- Hex Addr	0441	1089
x"00",	-- Hex Addr	0442	1090
x"00",	-- Hex Addr	0443	1091
x"00",	-- Hex Addr	0444	1092
x"00",	-- Hex Addr	0445	1093
x"00",	-- Hex Addr	0446	1094
x"00",	-- Hex Addr	0447	1095
x"00",	-- Hex Addr	0448	1096
x"00",	-- Hex Addr	0449	1097
x"00",	-- Hex Addr	044A	1098
x"00",	-- Hex Addr	044B	1099
x"00",	-- Hex Addr	044C	1100
x"00",	-- Hex Addr	044D	1101
x"00",	-- Hex Addr	044E	1102
x"00",	-- Hex Addr	044F	1103
x"00",	-- Hex Addr	0450	1104
x"00",	-- Hex Addr	0451	1105
x"00",	-- Hex Addr	0452	1106
x"00",	-- Hex Addr	0453	1107
x"00",	-- Hex Addr	0454	1108
x"00",	-- Hex Addr	0455	1109
x"00",	-- Hex Addr	0456	1110
x"00",	-- Hex Addr	0457	1111
x"00",	-- Hex Addr	0458	1112
x"00",	-- Hex Addr	0459	1113
x"00",	-- Hex Addr	045A	1114
x"00",	-- Hex Addr	045B	1115
x"00",	-- Hex Addr	045C	1116
x"00",	-- Hex Addr	045D	1117
x"00",	-- Hex Addr	045E	1118
x"00",	-- Hex Addr	045F	1119
x"00",	-- Hex Addr	0460	1120
x"00",	-- Hex Addr	0461	1121
x"00",	-- Hex Addr	0462	1122
x"00",	-- Hex Addr	0463	1123
x"00",	-- Hex Addr	0464	1124
x"00",	-- Hex Addr	0465	1125
x"00",	-- Hex Addr	0466	1126
x"00",	-- Hex Addr	0467	1127
x"00",	-- Hex Addr	0468	1128
x"00",	-- Hex Addr	0469	1129
x"00",	-- Hex Addr	046A	1130
x"00",	-- Hex Addr	046B	1131
x"00",	-- Hex Addr	046C	1132
x"00",	-- Hex Addr	046D	1133
x"00",	-- Hex Addr	046E	1134
x"00",	-- Hex Addr	046F	1135
x"00",	-- Hex Addr	0470	1136
x"00",	-- Hex Addr	0471	1137
x"00",	-- Hex Addr	0472	1138
x"00",	-- Hex Addr	0473	1139
x"00",	-- Hex Addr	0474	1140
x"00",	-- Hex Addr	0475	1141
x"00",	-- Hex Addr	0476	1142
x"00",	-- Hex Addr	0477	1143
x"00",	-- Hex Addr	0478	1144
x"00",	-- Hex Addr	0479	1145
x"00",	-- Hex Addr	047A	1146
x"00",	-- Hex Addr	047B	1147
x"00",	-- Hex Addr	047C	1148
x"00",	-- Hex Addr	047D	1149
x"00",	-- Hex Addr	047E	1150
x"00",	-- Hex Addr	047F	1151
x"00",	-- Hex Addr	0480	1152
x"00",	-- Hex Addr	0481	1153
x"00",	-- Hex Addr	0482	1154
x"00",	-- Hex Addr	0483	1155
x"00",	-- Hex Addr	0484	1156
x"00",	-- Hex Addr	0485	1157
x"00",	-- Hex Addr	0486	1158
x"00",	-- Hex Addr	0487	1159
x"00",	-- Hex Addr	0488	1160
x"00",	-- Hex Addr	0489	1161
x"00",	-- Hex Addr	048A	1162
x"00",	-- Hex Addr	048B	1163
x"00",	-- Hex Addr	048C	1164
x"00",	-- Hex Addr	048D	1165
x"00",	-- Hex Addr	048E	1166
x"00",	-- Hex Addr	048F	1167
x"00",	-- Hex Addr	0490	1168
x"00",	-- Hex Addr	0491	1169
x"00",	-- Hex Addr	0492	1170
x"00",	-- Hex Addr	0493	1171
x"00",	-- Hex Addr	0494	1172
x"00",	-- Hex Addr	0495	1173
x"00",	-- Hex Addr	0496	1174
x"00",	-- Hex Addr	0497	1175
x"00",	-- Hex Addr	0498	1176
x"00",	-- Hex Addr	0499	1177
x"00",	-- Hex Addr	049A	1178
x"00",	-- Hex Addr	049B	1179
x"00",	-- Hex Addr	049C	1180
x"00",	-- Hex Addr	049D	1181
x"00",	-- Hex Addr	049E	1182
x"00",	-- Hex Addr	049F	1183
x"00",	-- Hex Addr	04A0	1184
x"00",	-- Hex Addr	04A1	1185
x"00",	-- Hex Addr	04A2	1186
x"00",	-- Hex Addr	04A3	1187
x"00",	-- Hex Addr	04A4	1188
x"00",	-- Hex Addr	04A5	1189
x"00",	-- Hex Addr	04A6	1190
x"00",	-- Hex Addr	04A7	1191
x"00",	-- Hex Addr	04A8	1192
x"00",	-- Hex Addr	04A9	1193
x"00",	-- Hex Addr	04AA	1194
x"00",	-- Hex Addr	04AB	1195
x"00",	-- Hex Addr	04AC	1196
x"00",	-- Hex Addr	04AD	1197
x"00",	-- Hex Addr	04AE	1198
x"00",	-- Hex Addr	04AF	1199
x"00",	-- Hex Addr	04B0	1200
x"00",	-- Hex Addr	04B1	1201
x"00",	-- Hex Addr	04B2	1202
x"00",	-- Hex Addr	04B3	1203
x"00",	-- Hex Addr	04B4	1204
x"00",	-- Hex Addr	04B5	1205
x"00",	-- Hex Addr	04B6	1206
x"00",	-- Hex Addr	04B7	1207
x"00",	-- Hex Addr	04B8	1208
x"00",	-- Hex Addr	04B9	1209
x"00",	-- Hex Addr	04BA	1210
x"00",	-- Hex Addr	04BB	1211
x"00",	-- Hex Addr	04BC	1212
x"00",	-- Hex Addr	04BD	1213
x"00",	-- Hex Addr	04BE	1214
x"00",	-- Hex Addr	04BF	1215
x"00",	-- Hex Addr	04C0	1216
x"00",	-- Hex Addr	04C1	1217
x"00",	-- Hex Addr	04C2	1218
x"00",	-- Hex Addr	04C3	1219
x"00",	-- Hex Addr	04C4	1220
x"00",	-- Hex Addr	04C5	1221
x"00",	-- Hex Addr	04C6	1222
x"00",	-- Hex Addr	04C7	1223
x"00",	-- Hex Addr	04C8	1224
x"00",	-- Hex Addr	04C9	1225
x"00",	-- Hex Addr	04CA	1226
x"00",	-- Hex Addr	04CB	1227
x"00",	-- Hex Addr	04CC	1228
x"00",	-- Hex Addr	04CD	1229
x"00",	-- Hex Addr	04CE	1230
x"00",	-- Hex Addr	04CF	1231
x"00",	-- Hex Addr	04D0	1232
x"00",	-- Hex Addr	04D1	1233
x"00",	-- Hex Addr	04D2	1234
x"00",	-- Hex Addr	04D3	1235
x"00",	-- Hex Addr	04D4	1236
x"00",	-- Hex Addr	04D5	1237
x"00",	-- Hex Addr	04D6	1238
x"00",	-- Hex Addr	04D7	1239
x"00",	-- Hex Addr	04D8	1240
x"00",	-- Hex Addr	04D9	1241
x"00",	-- Hex Addr	04DA	1242
x"00",	-- Hex Addr	04DB	1243
x"00",	-- Hex Addr	04DC	1244
x"00",	-- Hex Addr	04DD	1245
x"00",	-- Hex Addr	04DE	1246
x"00",	-- Hex Addr	04DF	1247
x"00",	-- Hex Addr	04E0	1248
x"00",	-- Hex Addr	04E1	1249
x"00",	-- Hex Addr	04E2	1250
x"00",	-- Hex Addr	04E3	1251
x"00",	-- Hex Addr	04E4	1252
x"00",	-- Hex Addr	04E5	1253
x"00",	-- Hex Addr	04E6	1254
x"00",	-- Hex Addr	04E7	1255
x"00",	-- Hex Addr	04E8	1256
x"00",	-- Hex Addr	04E9	1257
x"00",	-- Hex Addr	04EA	1258
x"00",	-- Hex Addr	04EB	1259
x"00",	-- Hex Addr	04EC	1260
x"00",	-- Hex Addr	04ED	1261
x"00",	-- Hex Addr	04EE	1262
x"00",	-- Hex Addr	04EF	1263
x"00",	-- Hex Addr	04F0	1264
x"00",	-- Hex Addr	04F1	1265
x"00",	-- Hex Addr	04F2	1266
x"00",	-- Hex Addr	04F3	1267
x"00",	-- Hex Addr	04F4	1268
x"00",	-- Hex Addr	04F5	1269
x"00",	-- Hex Addr	04F6	1270
x"00",	-- Hex Addr	04F7	1271
x"00",	-- Hex Addr	04F8	1272
x"00",	-- Hex Addr	04F9	1273
x"00",	-- Hex Addr	04FA	1274
x"00",	-- Hex Addr	04FB	1275
x"00",	-- Hex Addr	04FC	1276
x"00",	-- Hex Addr	04FD	1277
x"00",	-- Hex Addr	04FE	1278
x"00",	-- Hex Addr	04FF	1279
x"00",	-- Hex Addr	0500	1280
x"00",	-- Hex Addr	0501	1281
x"00",	-- Hex Addr	0502	1282
x"00",	-- Hex Addr	0503	1283
x"00",	-- Hex Addr	0504	1284
x"00",	-- Hex Addr	0505	1285
x"00",	-- Hex Addr	0506	1286
x"00",	-- Hex Addr	0507	1287
x"00",	-- Hex Addr	0508	1288
x"00",	-- Hex Addr	0509	1289
x"00",	-- Hex Addr	050A	1290
x"00",	-- Hex Addr	050B	1291
x"00",	-- Hex Addr	050C	1292
x"00",	-- Hex Addr	050D	1293
x"00",	-- Hex Addr	050E	1294
x"00",	-- Hex Addr	050F	1295
x"00",	-- Hex Addr	0510	1296
x"00",	-- Hex Addr	0511	1297
x"00",	-- Hex Addr	0512	1298
x"00",	-- Hex Addr	0513	1299
x"00",	-- Hex Addr	0514	1300
x"00",	-- Hex Addr	0515	1301
x"00",	-- Hex Addr	0516	1302
x"00",	-- Hex Addr	0517	1303
x"00",	-- Hex Addr	0518	1304
x"00",	-- Hex Addr	0519	1305
x"00",	-- Hex Addr	051A	1306
x"00",	-- Hex Addr	051B	1307
x"00",	-- Hex Addr	051C	1308
x"00",	-- Hex Addr	051D	1309
x"00",	-- Hex Addr	051E	1310
x"00",	-- Hex Addr	051F	1311
x"00",	-- Hex Addr	0520	1312
x"00",	-- Hex Addr	0521	1313
x"00",	-- Hex Addr	0522	1314
x"00",	-- Hex Addr	0523	1315
x"00",	-- Hex Addr	0524	1316
x"00",	-- Hex Addr	0525	1317
x"00",	-- Hex Addr	0526	1318
x"00",	-- Hex Addr	0527	1319
x"00",	-- Hex Addr	0528	1320
x"00",	-- Hex Addr	0529	1321
x"00",	-- Hex Addr	052A	1322
x"00",	-- Hex Addr	052B	1323
x"00",	-- Hex Addr	052C	1324
x"00",	-- Hex Addr	052D	1325
x"00",	-- Hex Addr	052E	1326
x"00",	-- Hex Addr	052F	1327
x"00",	-- Hex Addr	0530	1328
x"00",	-- Hex Addr	0531	1329
x"00",	-- Hex Addr	0532	1330
x"00",	-- Hex Addr	0533	1331
x"00",	-- Hex Addr	0534	1332
x"00",	-- Hex Addr	0535	1333
x"00",	-- Hex Addr	0536	1334
x"00",	-- Hex Addr	0537	1335
x"00",	-- Hex Addr	0538	1336
x"00",	-- Hex Addr	0539	1337
x"00",	-- Hex Addr	053A	1338
x"00",	-- Hex Addr	053B	1339
x"00",	-- Hex Addr	053C	1340
x"00",	-- Hex Addr	053D	1341
x"00",	-- Hex Addr	053E	1342
x"00",	-- Hex Addr	053F	1343
x"00",	-- Hex Addr	0540	1344
x"00",	-- Hex Addr	0541	1345
x"00",	-- Hex Addr	0542	1346
x"00",	-- Hex Addr	0543	1347
x"00",	-- Hex Addr	0544	1348
x"00",	-- Hex Addr	0545	1349
x"00",	-- Hex Addr	0546	1350
x"00",	-- Hex Addr	0547	1351
x"00",	-- Hex Addr	0548	1352
x"00",	-- Hex Addr	0549	1353
x"00",	-- Hex Addr	054A	1354
x"00",	-- Hex Addr	054B	1355
x"00",	-- Hex Addr	054C	1356
x"00",	-- Hex Addr	054D	1357
x"00",	-- Hex Addr	054E	1358
x"00",	-- Hex Addr	054F	1359
x"00",	-- Hex Addr	0550	1360
x"00",	-- Hex Addr	0551	1361
x"00",	-- Hex Addr	0552	1362
x"00",	-- Hex Addr	0553	1363
x"00",	-- Hex Addr	0554	1364
x"00",	-- Hex Addr	0555	1365
x"00",	-- Hex Addr	0556	1366
x"00",	-- Hex Addr	0557	1367
x"00",	-- Hex Addr	0558	1368
x"00",	-- Hex Addr	0559	1369
x"00",	-- Hex Addr	055A	1370
x"00",	-- Hex Addr	055B	1371
x"00",	-- Hex Addr	055C	1372
x"00",	-- Hex Addr	055D	1373
x"00",	-- Hex Addr	055E	1374
x"00",	-- Hex Addr	055F	1375
x"00",	-- Hex Addr	0560	1376
x"00",	-- Hex Addr	0561	1377
x"00",	-- Hex Addr	0562	1378
x"00",	-- Hex Addr	0563	1379
x"00",	-- Hex Addr	0564	1380
x"00",	-- Hex Addr	0565	1381
x"00",	-- Hex Addr	0566	1382
x"00",	-- Hex Addr	0567	1383
x"00",	-- Hex Addr	0568	1384
x"00",	-- Hex Addr	0569	1385
x"00",	-- Hex Addr	056A	1386
x"00",	-- Hex Addr	056B	1387
x"00",	-- Hex Addr	056C	1388
x"00",	-- Hex Addr	056D	1389
x"00",	-- Hex Addr	056E	1390
x"00",	-- Hex Addr	056F	1391
x"00",	-- Hex Addr	0570	1392
x"00",	-- Hex Addr	0571	1393
x"00",	-- Hex Addr	0572	1394
x"00",	-- Hex Addr	0573	1395
x"00",	-- Hex Addr	0574	1396
x"00",	-- Hex Addr	0575	1397
x"00",	-- Hex Addr	0576	1398
x"00",	-- Hex Addr	0577	1399
x"00",	-- Hex Addr	0578	1400
x"00",	-- Hex Addr	0579	1401
x"00",	-- Hex Addr	057A	1402
x"00",	-- Hex Addr	057B	1403
x"00",	-- Hex Addr	057C	1404
x"00",	-- Hex Addr	057D	1405
x"00",	-- Hex Addr	057E	1406
x"00",	-- Hex Addr	057F	1407
x"00",	-- Hex Addr	0580	1408
x"00",	-- Hex Addr	0581	1409
x"00",	-- Hex Addr	0582	1410
x"00",	-- Hex Addr	0583	1411
x"00",	-- Hex Addr	0584	1412
x"00",	-- Hex Addr	0585	1413
x"00",	-- Hex Addr	0586	1414
x"00",	-- Hex Addr	0587	1415
x"00",	-- Hex Addr	0588	1416
x"00",	-- Hex Addr	0589	1417
x"00",	-- Hex Addr	058A	1418
x"00",	-- Hex Addr	058B	1419
x"00",	-- Hex Addr	058C	1420
x"00",	-- Hex Addr	058D	1421
x"00",	-- Hex Addr	058E	1422
x"00",	-- Hex Addr	058F	1423
x"00",	-- Hex Addr	0590	1424
x"00",	-- Hex Addr	0591	1425
x"00",	-- Hex Addr	0592	1426
x"00",	-- Hex Addr	0593	1427
x"00",	-- Hex Addr	0594	1428
x"00",	-- Hex Addr	0595	1429
x"00",	-- Hex Addr	0596	1430
x"00",	-- Hex Addr	0597	1431
x"00",	-- Hex Addr	0598	1432
x"00",	-- Hex Addr	0599	1433
x"00",	-- Hex Addr	059A	1434
x"00",	-- Hex Addr	059B	1435
x"00",	-- Hex Addr	059C	1436
x"00",	-- Hex Addr	059D	1437
x"00",	-- Hex Addr	059E	1438
x"00",	-- Hex Addr	059F	1439
x"00",	-- Hex Addr	05A0	1440
x"00",	-- Hex Addr	05A1	1441
x"00",	-- Hex Addr	05A2	1442
x"00",	-- Hex Addr	05A3	1443
x"00",	-- Hex Addr	05A4	1444
x"00",	-- Hex Addr	05A5	1445
x"00",	-- Hex Addr	05A6	1446
x"00",	-- Hex Addr	05A7	1447
x"00",	-- Hex Addr	05A8	1448
x"00",	-- Hex Addr	05A9	1449
x"00",	-- Hex Addr	05AA	1450
x"00",	-- Hex Addr	05AB	1451
x"00",	-- Hex Addr	05AC	1452
x"00",	-- Hex Addr	05AD	1453
x"00",	-- Hex Addr	05AE	1454
x"00",	-- Hex Addr	05AF	1455
x"00",	-- Hex Addr	05B0	1456
x"00",	-- Hex Addr	05B1	1457
x"00",	-- Hex Addr	05B2	1458
x"00",	-- Hex Addr	05B3	1459
x"00",	-- Hex Addr	05B4	1460
x"00",	-- Hex Addr	05B5	1461
x"00",	-- Hex Addr	05B6	1462
x"00",	-- Hex Addr	05B7	1463
x"00",	-- Hex Addr	05B8	1464
x"00",	-- Hex Addr	05B9	1465
x"00",	-- Hex Addr	05BA	1466
x"00",	-- Hex Addr	05BB	1467
x"00",	-- Hex Addr	05BC	1468
x"00",	-- Hex Addr	05BD	1469
x"00",	-- Hex Addr	05BE	1470
x"00",	-- Hex Addr	05BF	1471
x"00",	-- Hex Addr	05C0	1472
x"00",	-- Hex Addr	05C1	1473
x"00",	-- Hex Addr	05C2	1474
x"00",	-- Hex Addr	05C3	1475
x"00",	-- Hex Addr	05C4	1476
x"00",	-- Hex Addr	05C5	1477
x"00",	-- Hex Addr	05C6	1478
x"00",	-- Hex Addr	05C7	1479
x"00",	-- Hex Addr	05C8	1480
x"00",	-- Hex Addr	05C9	1481
x"00",	-- Hex Addr	05CA	1482
x"00",	-- Hex Addr	05CB	1483
x"00",	-- Hex Addr	05CC	1484
x"00",	-- Hex Addr	05CD	1485
x"00",	-- Hex Addr	05CE	1486
x"00",	-- Hex Addr	05CF	1487
x"00",	-- Hex Addr	05D0	1488
x"00",	-- Hex Addr	05D1	1489
x"00",	-- Hex Addr	05D2	1490
x"00",	-- Hex Addr	05D3	1491
x"00",	-- Hex Addr	05D4	1492
x"00",	-- Hex Addr	05D5	1493
x"00",	-- Hex Addr	05D6	1494
x"00",	-- Hex Addr	05D7	1495
x"00",	-- Hex Addr	05D8	1496
x"00",	-- Hex Addr	05D9	1497
x"00",	-- Hex Addr	05DA	1498
x"00",	-- Hex Addr	05DB	1499
x"00",	-- Hex Addr	05DC	1500
x"00",	-- Hex Addr	05DD	1501
x"00",	-- Hex Addr	05DE	1502
x"00",	-- Hex Addr	05DF	1503
x"00",	-- Hex Addr	05E0	1504
x"00",	-- Hex Addr	05E1	1505
x"00",	-- Hex Addr	05E2	1506
x"00",	-- Hex Addr	05E3	1507
x"00",	-- Hex Addr	05E4	1508
x"00",	-- Hex Addr	05E5	1509
x"00",	-- Hex Addr	05E6	1510
x"00",	-- Hex Addr	05E7	1511
x"00",	-- Hex Addr	05E8	1512
x"00",	-- Hex Addr	05E9	1513
x"00",	-- Hex Addr	05EA	1514
x"00",	-- Hex Addr	05EB	1515
x"00",	-- Hex Addr	05EC	1516
x"00",	-- Hex Addr	05ED	1517
x"00",	-- Hex Addr	05EE	1518
x"00",	-- Hex Addr	05EF	1519
x"00",	-- Hex Addr	05F0	1520
x"00",	-- Hex Addr	05F1	1521
x"00",	-- Hex Addr	05F2	1522
x"00",	-- Hex Addr	05F3	1523
x"00",	-- Hex Addr	05F4	1524
x"00",	-- Hex Addr	05F5	1525
x"00",	-- Hex Addr	05F6	1526
x"00",	-- Hex Addr	05F7	1527
x"00",	-- Hex Addr	05F8	1528
x"00",	-- Hex Addr	05F9	1529
x"00",	-- Hex Addr	05FA	1530
x"00",	-- Hex Addr	05FB	1531
x"00",	-- Hex Addr	05FC	1532
x"00",	-- Hex Addr	05FD	1533
x"00",	-- Hex Addr	05FE	1534
x"00",	-- Hex Addr	05FF	1535
x"00",	-- Hex Addr	0600	1536
x"00",	-- Hex Addr	0601	1537
x"00",	-- Hex Addr	0602	1538
x"00",	-- Hex Addr	0603	1539
x"00",	-- Hex Addr	0604	1540
x"00",	-- Hex Addr	0605	1541
x"00",	-- Hex Addr	0606	1542
x"00",	-- Hex Addr	0607	1543
x"00",	-- Hex Addr	0608	1544
x"00",	-- Hex Addr	0609	1545
x"00",	-- Hex Addr	060A	1546
x"00",	-- Hex Addr	060B	1547
x"00",	-- Hex Addr	060C	1548
x"00",	-- Hex Addr	060D	1549
x"00",	-- Hex Addr	060E	1550
x"00",	-- Hex Addr	060F	1551
x"00",	-- Hex Addr	0610	1552
x"00",	-- Hex Addr	0611	1553
x"00",	-- Hex Addr	0612	1554
x"00",	-- Hex Addr	0613	1555
x"00",	-- Hex Addr	0614	1556
x"00",	-- Hex Addr	0615	1557
x"00",	-- Hex Addr	0616	1558
x"00",	-- Hex Addr	0617	1559
x"00",	-- Hex Addr	0618	1560
x"00",	-- Hex Addr	0619	1561
x"00",	-- Hex Addr	061A	1562
x"00",	-- Hex Addr	061B	1563
x"00",	-- Hex Addr	061C	1564
x"00",	-- Hex Addr	061D	1565
x"00",	-- Hex Addr	061E	1566
x"00",	-- Hex Addr	061F	1567
x"00",	-- Hex Addr	0620	1568
x"00",	-- Hex Addr	0621	1569
x"00",	-- Hex Addr	0622	1570
x"00",	-- Hex Addr	0623	1571
x"00",	-- Hex Addr	0624	1572
x"00",	-- Hex Addr	0625	1573
x"00",	-- Hex Addr	0626	1574
x"00",	-- Hex Addr	0627	1575
x"00",	-- Hex Addr	0628	1576
x"00",	-- Hex Addr	0629	1577
x"00",	-- Hex Addr	062A	1578
x"00",	-- Hex Addr	062B	1579
x"00",	-- Hex Addr	062C	1580
x"00",	-- Hex Addr	062D	1581
x"00",	-- Hex Addr	062E	1582
x"00",	-- Hex Addr	062F	1583
x"00",	-- Hex Addr	0630	1584
x"00",	-- Hex Addr	0631	1585
x"00",	-- Hex Addr	0632	1586
x"00",	-- Hex Addr	0633	1587
x"00",	-- Hex Addr	0634	1588
x"00",	-- Hex Addr	0635	1589
x"00",	-- Hex Addr	0636	1590
x"00",	-- Hex Addr	0637	1591
x"00",	-- Hex Addr	0638	1592
x"00",	-- Hex Addr	0639	1593
x"00",	-- Hex Addr	063A	1594
x"00",	-- Hex Addr	063B	1595
x"00",	-- Hex Addr	063C	1596
x"00",	-- Hex Addr	063D	1597
x"00",	-- Hex Addr	063E	1598
x"00",	-- Hex Addr	063F	1599
x"00",	-- Hex Addr	0640	1600
x"00",	-- Hex Addr	0641	1601
x"00",	-- Hex Addr	0642	1602
x"00",	-- Hex Addr	0643	1603
x"00",	-- Hex Addr	0644	1604
x"00",	-- Hex Addr	0645	1605
x"00",	-- Hex Addr	0646	1606
x"00",	-- Hex Addr	0647	1607
x"00",	-- Hex Addr	0648	1608
x"00",	-- Hex Addr	0649	1609
x"00",	-- Hex Addr	064A	1610
x"00",	-- Hex Addr	064B	1611
x"00",	-- Hex Addr	064C	1612
x"00",	-- Hex Addr	064D	1613
x"00",	-- Hex Addr	064E	1614
x"00",	-- Hex Addr	064F	1615
x"00",	-- Hex Addr	0650	1616
x"00",	-- Hex Addr	0651	1617
x"00",	-- Hex Addr	0652	1618
x"00",	-- Hex Addr	0653	1619
x"00",	-- Hex Addr	0654	1620
x"00",	-- Hex Addr	0655	1621
x"00",	-- Hex Addr	0656	1622
x"00",	-- Hex Addr	0657	1623
x"00",	-- Hex Addr	0658	1624
x"00",	-- Hex Addr	0659	1625
x"00",	-- Hex Addr	065A	1626
x"00",	-- Hex Addr	065B	1627
x"00",	-- Hex Addr	065C	1628
x"00",	-- Hex Addr	065D	1629
x"00",	-- Hex Addr	065E	1630
x"00",	-- Hex Addr	065F	1631
x"00",	-- Hex Addr	0660	1632
x"00",	-- Hex Addr	0661	1633
x"00",	-- Hex Addr	0662	1634
x"00",	-- Hex Addr	0663	1635
x"00",	-- Hex Addr	0664	1636
x"00",	-- Hex Addr	0665	1637
x"00",	-- Hex Addr	0666	1638
x"00",	-- Hex Addr	0667	1639
x"00",	-- Hex Addr	0668	1640
x"00",	-- Hex Addr	0669	1641
x"00",	-- Hex Addr	066A	1642
x"00",	-- Hex Addr	066B	1643
x"00",	-- Hex Addr	066C	1644
x"00",	-- Hex Addr	066D	1645
x"00",	-- Hex Addr	066E	1646
x"00",	-- Hex Addr	066F	1647
x"00",	-- Hex Addr	0670	1648
x"00",	-- Hex Addr	0671	1649
x"00",	-- Hex Addr	0672	1650
x"00",	-- Hex Addr	0673	1651
x"00",	-- Hex Addr	0674	1652
x"00",	-- Hex Addr	0675	1653
x"00",	-- Hex Addr	0676	1654
x"00",	-- Hex Addr	0677	1655
x"00",	-- Hex Addr	0678	1656
x"00",	-- Hex Addr	0679	1657
x"00",	-- Hex Addr	067A	1658
x"00",	-- Hex Addr	067B	1659
x"00",	-- Hex Addr	067C	1660
x"00",	-- Hex Addr	067D	1661
x"00",	-- Hex Addr	067E	1662
x"00",	-- Hex Addr	067F	1663
x"00",	-- Hex Addr	0680	1664
x"00",	-- Hex Addr	0681	1665
x"00",	-- Hex Addr	0682	1666
x"00",	-- Hex Addr	0683	1667
x"00",	-- Hex Addr	0684	1668
x"00",	-- Hex Addr	0685	1669
x"00",	-- Hex Addr	0686	1670
x"00",	-- Hex Addr	0687	1671
x"00",	-- Hex Addr	0688	1672
x"00",	-- Hex Addr	0689	1673
x"00",	-- Hex Addr	068A	1674
x"00",	-- Hex Addr	068B	1675
x"00",	-- Hex Addr	068C	1676
x"00",	-- Hex Addr	068D	1677
x"00",	-- Hex Addr	068E	1678
x"00",	-- Hex Addr	068F	1679
x"00",	-- Hex Addr	0690	1680
x"00",	-- Hex Addr	0691	1681
x"00",	-- Hex Addr	0692	1682
x"00",	-- Hex Addr	0693	1683
x"00",	-- Hex Addr	0694	1684
x"00",	-- Hex Addr	0695	1685
x"00",	-- Hex Addr	0696	1686
x"00",	-- Hex Addr	0697	1687
x"00",	-- Hex Addr	0698	1688
x"00",	-- Hex Addr	0699	1689
x"00",	-- Hex Addr	069A	1690
x"00",	-- Hex Addr	069B	1691
x"00",	-- Hex Addr	069C	1692
x"00",	-- Hex Addr	069D	1693
x"00",	-- Hex Addr	069E	1694
x"00",	-- Hex Addr	069F	1695
x"00",	-- Hex Addr	06A0	1696
x"00",	-- Hex Addr	06A1	1697
x"00",	-- Hex Addr	06A2	1698
x"00",	-- Hex Addr	06A3	1699
x"00",	-- Hex Addr	06A4	1700
x"00",	-- Hex Addr	06A5	1701
x"00",	-- Hex Addr	06A6	1702
x"00",	-- Hex Addr	06A7	1703
x"00",	-- Hex Addr	06A8	1704
x"00",	-- Hex Addr	06A9	1705
x"00",	-- Hex Addr	06AA	1706
x"00",	-- Hex Addr	06AB	1707
x"00",	-- Hex Addr	06AC	1708
x"00",	-- Hex Addr	06AD	1709
x"00",	-- Hex Addr	06AE	1710
x"00",	-- Hex Addr	06AF	1711
x"00",	-- Hex Addr	06B0	1712
x"00",	-- Hex Addr	06B1	1713
x"00",	-- Hex Addr	06B2	1714
x"00",	-- Hex Addr	06B3	1715
x"00",	-- Hex Addr	06B4	1716
x"00",	-- Hex Addr	06B5	1717
x"00",	-- Hex Addr	06B6	1718
x"00",	-- Hex Addr	06B7	1719
x"00",	-- Hex Addr	06B8	1720
x"00",	-- Hex Addr	06B9	1721
x"00",	-- Hex Addr	06BA	1722
x"00",	-- Hex Addr	06BB	1723
x"00",	-- Hex Addr	06BC	1724
x"00",	-- Hex Addr	06BD	1725
x"00",	-- Hex Addr	06BE	1726
x"00",	-- Hex Addr	06BF	1727
x"00",	-- Hex Addr	06C0	1728
x"00",	-- Hex Addr	06C1	1729
x"00",	-- Hex Addr	06C2	1730
x"00",	-- Hex Addr	06C3	1731
x"00",	-- Hex Addr	06C4	1732
x"00",	-- Hex Addr	06C5	1733
x"00",	-- Hex Addr	06C6	1734
x"00",	-- Hex Addr	06C7	1735
x"00",	-- Hex Addr	06C8	1736
x"00",	-- Hex Addr	06C9	1737
x"00",	-- Hex Addr	06CA	1738
x"00",	-- Hex Addr	06CB	1739
x"00",	-- Hex Addr	06CC	1740
x"00",	-- Hex Addr	06CD	1741
x"00",	-- Hex Addr	06CE	1742
x"00",	-- Hex Addr	06CF	1743
x"00",	-- Hex Addr	06D0	1744
x"00",	-- Hex Addr	06D1	1745
x"00",	-- Hex Addr	06D2	1746
x"00",	-- Hex Addr	06D3	1747
x"00",	-- Hex Addr	06D4	1748
x"00",	-- Hex Addr	06D5	1749
x"00",	-- Hex Addr	06D6	1750
x"00",	-- Hex Addr	06D7	1751
x"00",	-- Hex Addr	06D8	1752
x"00",	-- Hex Addr	06D9	1753
x"00",	-- Hex Addr	06DA	1754
x"00",	-- Hex Addr	06DB	1755
x"00",	-- Hex Addr	06DC	1756
x"00",	-- Hex Addr	06DD	1757
x"00",	-- Hex Addr	06DE	1758
x"00",	-- Hex Addr	06DF	1759
x"00",	-- Hex Addr	06E0	1760
x"00",	-- Hex Addr	06E1	1761
x"00",	-- Hex Addr	06E2	1762
x"00",	-- Hex Addr	06E3	1763
x"00",	-- Hex Addr	06E4	1764
x"00",	-- Hex Addr	06E5	1765
x"00",	-- Hex Addr	06E6	1766
x"00",	-- Hex Addr	06E7	1767
x"00",	-- Hex Addr	06E8	1768
x"00",	-- Hex Addr	06E9	1769
x"00",	-- Hex Addr	06EA	1770
x"00",	-- Hex Addr	06EB	1771
x"00",	-- Hex Addr	06EC	1772
x"00",	-- Hex Addr	06ED	1773
x"00",	-- Hex Addr	06EE	1774
x"00",	-- Hex Addr	06EF	1775
x"00",	-- Hex Addr	06F0	1776
x"00",	-- Hex Addr	06F1	1777
x"00",	-- Hex Addr	06F2	1778
x"00",	-- Hex Addr	06F3	1779
x"00",	-- Hex Addr	06F4	1780
x"00",	-- Hex Addr	06F5	1781
x"00",	-- Hex Addr	06F6	1782
x"00",	-- Hex Addr	06F7	1783
x"00",	-- Hex Addr	06F8	1784
x"00",	-- Hex Addr	06F9	1785
x"00",	-- Hex Addr	06FA	1786
x"00",	-- Hex Addr	06FB	1787
x"00",	-- Hex Addr	06FC	1788
x"00",	-- Hex Addr	06FD	1789
x"00",	-- Hex Addr	06FE	1790
x"00",	-- Hex Addr	06FF	1791
x"00",	-- Hex Addr	0700	1792
x"00",	-- Hex Addr	0701	1793
x"00",	-- Hex Addr	0702	1794
x"00",	-- Hex Addr	0703	1795
x"00",	-- Hex Addr	0704	1796
x"00",	-- Hex Addr	0705	1797
x"00",	-- Hex Addr	0706	1798
x"00",	-- Hex Addr	0707	1799
x"00",	-- Hex Addr	0708	1800
x"00",	-- Hex Addr	0709	1801
x"00",	-- Hex Addr	070A	1802
x"00",	-- Hex Addr	070B	1803
x"00",	-- Hex Addr	070C	1804
x"00",	-- Hex Addr	070D	1805
x"00",	-- Hex Addr	070E	1806
x"00",	-- Hex Addr	070F	1807
x"00",	-- Hex Addr	0710	1808
x"00",	-- Hex Addr	0711	1809
x"00",	-- Hex Addr	0712	1810
x"00",	-- Hex Addr	0713	1811
x"00",	-- Hex Addr	0714	1812
x"00",	-- Hex Addr	0715	1813
x"00",	-- Hex Addr	0716	1814
x"00",	-- Hex Addr	0717	1815
x"00",	-- Hex Addr	0718	1816
x"00",	-- Hex Addr	0719	1817
x"00",	-- Hex Addr	071A	1818
x"00",	-- Hex Addr	071B	1819
x"00",	-- Hex Addr	071C	1820
x"00",	-- Hex Addr	071D	1821
x"00",	-- Hex Addr	071E	1822
x"00",	-- Hex Addr	071F	1823
x"00",	-- Hex Addr	0720	1824
x"00",	-- Hex Addr	0721	1825
x"00",	-- Hex Addr	0722	1826
x"00",	-- Hex Addr	0723	1827
x"00",	-- Hex Addr	0724	1828
x"00",	-- Hex Addr	0725	1829
x"00",	-- Hex Addr	0726	1830
x"00",	-- Hex Addr	0727	1831
x"00",	-- Hex Addr	0728	1832
x"00",	-- Hex Addr	0729	1833
x"00",	-- Hex Addr	072A	1834
x"00",	-- Hex Addr	072B	1835
x"00",	-- Hex Addr	072C	1836
x"00",	-- Hex Addr	072D	1837
x"00",	-- Hex Addr	072E	1838
x"00",	-- Hex Addr	072F	1839
x"00",	-- Hex Addr	0730	1840
x"00",	-- Hex Addr	0731	1841
x"00",	-- Hex Addr	0732	1842
x"00",	-- Hex Addr	0733	1843
x"00",	-- Hex Addr	0734	1844
x"00",	-- Hex Addr	0735	1845
x"00",	-- Hex Addr	0736	1846
x"00",	-- Hex Addr	0737	1847
x"00",	-- Hex Addr	0738	1848
x"00",	-- Hex Addr	0739	1849
x"00",	-- Hex Addr	073A	1850
x"00",	-- Hex Addr	073B	1851
x"00",	-- Hex Addr	073C	1852
x"00",	-- Hex Addr	073D	1853
x"00",	-- Hex Addr	073E	1854
x"00",	-- Hex Addr	073F	1855
x"00",	-- Hex Addr	0740	1856
x"00",	-- Hex Addr	0741	1857
x"00",	-- Hex Addr	0742	1858
x"00",	-- Hex Addr	0743	1859
x"00",	-- Hex Addr	0744	1860
x"00",	-- Hex Addr	0745	1861
x"00",	-- Hex Addr	0746	1862
x"00",	-- Hex Addr	0747	1863
x"00",	-- Hex Addr	0748	1864
x"00",	-- Hex Addr	0749	1865
x"00",	-- Hex Addr	074A	1866
x"00",	-- Hex Addr	074B	1867
x"00",	-- Hex Addr	074C	1868
x"00",	-- Hex Addr	074D	1869
x"00",	-- Hex Addr	074E	1870
x"00",	-- Hex Addr	074F	1871
x"00",	-- Hex Addr	0750	1872
x"00",	-- Hex Addr	0751	1873
x"00",	-- Hex Addr	0752	1874
x"00",	-- Hex Addr	0753	1875
x"00",	-- Hex Addr	0754	1876
x"00",	-- Hex Addr	0755	1877
x"00",	-- Hex Addr	0756	1878
x"00",	-- Hex Addr	0757	1879
x"00",	-- Hex Addr	0758	1880
x"00",	-- Hex Addr	0759	1881
x"00",	-- Hex Addr	075A	1882
x"00",	-- Hex Addr	075B	1883
x"00",	-- Hex Addr	075C	1884
x"00",	-- Hex Addr	075D	1885
x"00",	-- Hex Addr	075E	1886
x"00",	-- Hex Addr	075F	1887
x"00",	-- Hex Addr	0760	1888
x"00",	-- Hex Addr	0761	1889
x"00",	-- Hex Addr	0762	1890
x"00",	-- Hex Addr	0763	1891
x"00",	-- Hex Addr	0764	1892
x"00",	-- Hex Addr	0765	1893
x"00",	-- Hex Addr	0766	1894
x"00",	-- Hex Addr	0767	1895
x"00",	-- Hex Addr	0768	1896
x"00",	-- Hex Addr	0769	1897
x"00",	-- Hex Addr	076A	1898
x"00",	-- Hex Addr	076B	1899
x"00",	-- Hex Addr	076C	1900
x"00",	-- Hex Addr	076D	1901
x"00",	-- Hex Addr	076E	1902
x"00",	-- Hex Addr	076F	1903
x"00",	-- Hex Addr	0770	1904
x"00",	-- Hex Addr	0771	1905
x"00",	-- Hex Addr	0772	1906
x"00",	-- Hex Addr	0773	1907
x"00",	-- Hex Addr	0774	1908
x"00",	-- Hex Addr	0775	1909
x"00",	-- Hex Addr	0776	1910
x"00",	-- Hex Addr	0777	1911
x"00",	-- Hex Addr	0778	1912
x"00",	-- Hex Addr	0779	1913
x"00",	-- Hex Addr	077A	1914
x"00",	-- Hex Addr	077B	1915
x"00",	-- Hex Addr	077C	1916
x"00",	-- Hex Addr	077D	1917
x"00",	-- Hex Addr	077E	1918
x"00",	-- Hex Addr	077F	1919
x"00",	-- Hex Addr	0780	1920
x"00",	-- Hex Addr	0781	1921
x"00",	-- Hex Addr	0782	1922
x"00",	-- Hex Addr	0783	1923
x"00",	-- Hex Addr	0784	1924
x"00",	-- Hex Addr	0785	1925
x"00",	-- Hex Addr	0786	1926
x"00",	-- Hex Addr	0787	1927
x"00",	-- Hex Addr	0788	1928
x"00",	-- Hex Addr	0789	1929
x"00",	-- Hex Addr	078A	1930
x"00",	-- Hex Addr	078B	1931
x"00",	-- Hex Addr	078C	1932
x"00",	-- Hex Addr	078D	1933
x"00",	-- Hex Addr	078E	1934
x"00",	-- Hex Addr	078F	1935
x"00",	-- Hex Addr	0790	1936
x"00",	-- Hex Addr	0791	1937
x"00",	-- Hex Addr	0792	1938
x"00",	-- Hex Addr	0793	1939
x"00",	-- Hex Addr	0794	1940
x"00",	-- Hex Addr	0795	1941
x"00",	-- Hex Addr	0796	1942
x"00",	-- Hex Addr	0797	1943
x"00",	-- Hex Addr	0798	1944
x"00",	-- Hex Addr	0799	1945
x"00",	-- Hex Addr	079A	1946
x"00",	-- Hex Addr	079B	1947
x"00",	-- Hex Addr	079C	1948
x"00",	-- Hex Addr	079D	1949
x"00",	-- Hex Addr	079E	1950
x"00",	-- Hex Addr	079F	1951
x"00",	-- Hex Addr	07A0	1952
x"00",	-- Hex Addr	07A1	1953
x"00",	-- Hex Addr	07A2	1954
x"00",	-- Hex Addr	07A3	1955
x"00",	-- Hex Addr	07A4	1956
x"00",	-- Hex Addr	07A5	1957
x"00",	-- Hex Addr	07A6	1958
x"00",	-- Hex Addr	07A7	1959
x"00",	-- Hex Addr	07A8	1960
x"00",	-- Hex Addr	07A9	1961
x"00",	-- Hex Addr	07AA	1962
x"00",	-- Hex Addr	07AB	1963
x"00",	-- Hex Addr	07AC	1964
x"00",	-- Hex Addr	07AD	1965
x"00",	-- Hex Addr	07AE	1966
x"00",	-- Hex Addr	07AF	1967
x"00",	-- Hex Addr	07B0	1968
x"00",	-- Hex Addr	07B1	1969
x"00",	-- Hex Addr	07B2	1970
x"00",	-- Hex Addr	07B3	1971
x"00",	-- Hex Addr	07B4	1972
x"00",	-- Hex Addr	07B5	1973
x"00",	-- Hex Addr	07B6	1974
x"00",	-- Hex Addr	07B7	1975
x"00",	-- Hex Addr	07B8	1976
x"00",	-- Hex Addr	07B9	1977
x"00",	-- Hex Addr	07BA	1978
x"00",	-- Hex Addr	07BB	1979
x"00",	-- Hex Addr	07BC	1980
x"00",	-- Hex Addr	07BD	1981
x"00",	-- Hex Addr	07BE	1982
x"00",	-- Hex Addr	07BF	1983
x"00",	-- Hex Addr	07C0	1984
x"00",	-- Hex Addr	07C1	1985
x"00",	-- Hex Addr	07C2	1986
x"00",	-- Hex Addr	07C3	1987
x"00",	-- Hex Addr	07C4	1988
x"00",	-- Hex Addr	07C5	1989
x"00",	-- Hex Addr	07C6	1990
x"00",	-- Hex Addr	07C7	1991
x"00",	-- Hex Addr	07C8	1992
x"00",	-- Hex Addr	07C9	1993
x"00",	-- Hex Addr	07CA	1994
x"00",	-- Hex Addr	07CB	1995
x"00",	-- Hex Addr	07CC	1996
x"00",	-- Hex Addr	07CD	1997
x"00",	-- Hex Addr	07CE	1998
x"00",	-- Hex Addr	07CF	1999
x"00",	-- Hex Addr	07D0	2000
x"00",	-- Hex Addr	07D1	2001
x"00",	-- Hex Addr	07D2	2002
x"00",	-- Hex Addr	07D3	2003
x"00",	-- Hex Addr	07D4	2004
x"00",	-- Hex Addr	07D5	2005
x"00",	-- Hex Addr	07D6	2006
x"00",	-- Hex Addr	07D7	2007
x"00",	-- Hex Addr	07D8	2008
x"00",	-- Hex Addr	07D9	2009
x"00",	-- Hex Addr	07DA	2010
x"00",	-- Hex Addr	07DB	2011
x"00",	-- Hex Addr	07DC	2012
x"00",	-- Hex Addr	07DD	2013
x"00",	-- Hex Addr	07DE	2014
x"00",	-- Hex Addr	07DF	2015
x"00",	-- Hex Addr	07E0	2016
x"00",	-- Hex Addr	07E1	2017
x"00",	-- Hex Addr	07E2	2018
x"00",	-- Hex Addr	07E3	2019
x"00",	-- Hex Addr	07E4	2020
x"00",	-- Hex Addr	07E5	2021
x"00",	-- Hex Addr	07E6	2022
x"00",	-- Hex Addr	07E7	2023
x"00",	-- Hex Addr	07E8	2024
x"00",	-- Hex Addr	07E9	2025
x"00",	-- Hex Addr	07EA	2026
x"00",	-- Hex Addr	07EB	2027
x"00",	-- Hex Addr	07EC	2028
x"00",	-- Hex Addr	07ED	2029
x"00",	-- Hex Addr	07EE	2030
x"00",	-- Hex Addr	07EF	2031
x"00",	-- Hex Addr	07F0	2032
x"00",	-- Hex Addr	07F1	2033
x"00",	-- Hex Addr	07F2	2034
x"00",	-- Hex Addr	07F3	2035
x"00",	-- Hex Addr	07F4	2036
x"00",	-- Hex Addr	07F5	2037
x"00",	-- Hex Addr	07F6	2038
x"00",	-- Hex Addr	07F7	2039
x"00",	-- Hex Addr	07F8	2040
x"00",	-- Hex Addr	07F9	2041
x"00",	-- Hex Addr	07FA	2042
x"00",	-- Hex Addr	07FB	2043
x"00",	-- Hex Addr	07FC	2044
x"00",	-- Hex Addr	07FD	2045
x"00",	-- Hex Addr	07FE	2046
x"00",	-- Hex Addr	07FF	2047
x"00",	-- Hex Addr	0800	2048
x"00",	-- Hex Addr	0801	2049
x"00",	-- Hex Addr	0802	2050
x"00",	-- Hex Addr	0803	2051
x"00",	-- Hex Addr	0804	2052
x"00",	-- Hex Addr	0805	2053
x"00",	-- Hex Addr	0806	2054
x"00",	-- Hex Addr	0807	2055
x"00",	-- Hex Addr	0808	2056
x"00",	-- Hex Addr	0809	2057
x"00",	-- Hex Addr	080A	2058
x"00",	-- Hex Addr	080B	2059
x"00",	-- Hex Addr	080C	2060
x"00",	-- Hex Addr	080D	2061
x"00",	-- Hex Addr	080E	2062
x"00",	-- Hex Addr	080F	2063
x"00",	-- Hex Addr	0810	2064
x"00",	-- Hex Addr	0811	2065
x"00",	-- Hex Addr	0812	2066
x"00",	-- Hex Addr	0813	2067
x"00",	-- Hex Addr	0814	2068
x"00",	-- Hex Addr	0815	2069
x"00",	-- Hex Addr	0816	2070
x"00",	-- Hex Addr	0817	2071
x"00",	-- Hex Addr	0818	2072
x"00",	-- Hex Addr	0819	2073
x"00",	-- Hex Addr	081A	2074
x"00",	-- Hex Addr	081B	2075
x"00",	-- Hex Addr	081C	2076
x"00",	-- Hex Addr	081D	2077
x"00",	-- Hex Addr	081E	2078
x"00",	-- Hex Addr	081F	2079
x"00",	-- Hex Addr	0820	2080
x"00",	-- Hex Addr	0821	2081
x"00",	-- Hex Addr	0822	2082
x"00",	-- Hex Addr	0823	2083
x"00",	-- Hex Addr	0824	2084
x"00",	-- Hex Addr	0825	2085
x"00",	-- Hex Addr	0826	2086
x"00",	-- Hex Addr	0827	2087
x"00",	-- Hex Addr	0828	2088
x"00",	-- Hex Addr	0829	2089
x"00",	-- Hex Addr	082A	2090
x"00",	-- Hex Addr	082B	2091
x"00",	-- Hex Addr	082C	2092
x"00",	-- Hex Addr	082D	2093
x"00",	-- Hex Addr	082E	2094
x"00",	-- Hex Addr	082F	2095
x"00",	-- Hex Addr	0830	2096
x"00",	-- Hex Addr	0831	2097
x"00",	-- Hex Addr	0832	2098
x"00",	-- Hex Addr	0833	2099
x"00",	-- Hex Addr	0834	2100
x"00",	-- Hex Addr	0835	2101
x"00",	-- Hex Addr	0836	2102
x"00",	-- Hex Addr	0837	2103
x"00",	-- Hex Addr	0838	2104
x"00",	-- Hex Addr	0839	2105
x"00",	-- Hex Addr	083A	2106
x"00",	-- Hex Addr	083B	2107
x"00",	-- Hex Addr	083C	2108
x"00",	-- Hex Addr	083D	2109
x"00",	-- Hex Addr	083E	2110
x"00",	-- Hex Addr	083F	2111
x"00",	-- Hex Addr	0840	2112
x"00",	-- Hex Addr	0841	2113
x"00",	-- Hex Addr	0842	2114
x"00",	-- Hex Addr	0843	2115
x"00",	-- Hex Addr	0844	2116
x"00",	-- Hex Addr	0845	2117
x"00",	-- Hex Addr	0846	2118
x"00",	-- Hex Addr	0847	2119
x"00",	-- Hex Addr	0848	2120
x"00",	-- Hex Addr	0849	2121
x"00",	-- Hex Addr	084A	2122
x"00",	-- Hex Addr	084B	2123
x"00",	-- Hex Addr	084C	2124
x"00",	-- Hex Addr	084D	2125
x"00",	-- Hex Addr	084E	2126
x"00",	-- Hex Addr	084F	2127
x"00",	-- Hex Addr	0850	2128
x"00",	-- Hex Addr	0851	2129
x"00",	-- Hex Addr	0852	2130
x"00",	-- Hex Addr	0853	2131
x"00",	-- Hex Addr	0854	2132
x"00",	-- Hex Addr	0855	2133
x"00",	-- Hex Addr	0856	2134
x"00",	-- Hex Addr	0857	2135
x"00",	-- Hex Addr	0858	2136
x"00",	-- Hex Addr	0859	2137
x"00",	-- Hex Addr	085A	2138
x"00",	-- Hex Addr	085B	2139
x"00",	-- Hex Addr	085C	2140
x"00",	-- Hex Addr	085D	2141
x"00",	-- Hex Addr	085E	2142
x"00",	-- Hex Addr	085F	2143
x"00",	-- Hex Addr	0860	2144
x"00",	-- Hex Addr	0861	2145
x"00",	-- Hex Addr	0862	2146
x"00",	-- Hex Addr	0863	2147
x"00",	-- Hex Addr	0864	2148
x"00",	-- Hex Addr	0865	2149
x"00",	-- Hex Addr	0866	2150
x"00",	-- Hex Addr	0867	2151
x"00",	-- Hex Addr	0868	2152
x"00",	-- Hex Addr	0869	2153
x"00",	-- Hex Addr	086A	2154
x"00",	-- Hex Addr	086B	2155
x"00",	-- Hex Addr	086C	2156
x"00",	-- Hex Addr	086D	2157
x"00",	-- Hex Addr	086E	2158
x"00",	-- Hex Addr	086F	2159
x"00",	-- Hex Addr	0870	2160
x"00",	-- Hex Addr	0871	2161
x"00",	-- Hex Addr	0872	2162
x"00",	-- Hex Addr	0873	2163
x"00",	-- Hex Addr	0874	2164
x"00",	-- Hex Addr	0875	2165
x"00",	-- Hex Addr	0876	2166
x"00",	-- Hex Addr	0877	2167
x"00",	-- Hex Addr	0878	2168
x"00",	-- Hex Addr	0879	2169
x"00",	-- Hex Addr	087A	2170
x"00",	-- Hex Addr	087B	2171
x"00",	-- Hex Addr	087C	2172
x"00",	-- Hex Addr	087D	2173
x"00",	-- Hex Addr	087E	2174
x"00",	-- Hex Addr	087F	2175
x"00",	-- Hex Addr	0880	2176
x"00",	-- Hex Addr	0881	2177
x"00",	-- Hex Addr	0882	2178
x"00",	-- Hex Addr	0883	2179
x"00",	-- Hex Addr	0884	2180
x"00",	-- Hex Addr	0885	2181
x"00",	-- Hex Addr	0886	2182
x"00",	-- Hex Addr	0887	2183
x"00",	-- Hex Addr	0888	2184
x"00",	-- Hex Addr	0889	2185
x"00",	-- Hex Addr	088A	2186
x"00",	-- Hex Addr	088B	2187
x"00",	-- Hex Addr	088C	2188
x"00",	-- Hex Addr	088D	2189
x"00",	-- Hex Addr	088E	2190
x"00",	-- Hex Addr	088F	2191
x"00",	-- Hex Addr	0890	2192
x"00",	-- Hex Addr	0891	2193
x"00",	-- Hex Addr	0892	2194
x"00",	-- Hex Addr	0893	2195
x"00",	-- Hex Addr	0894	2196
x"00",	-- Hex Addr	0895	2197
x"00",	-- Hex Addr	0896	2198
x"00",	-- Hex Addr	0897	2199
x"00",	-- Hex Addr	0898	2200
x"00",	-- Hex Addr	0899	2201
x"00",	-- Hex Addr	089A	2202
x"00",	-- Hex Addr	089B	2203
x"00",	-- Hex Addr	089C	2204
x"00",	-- Hex Addr	089D	2205
x"00",	-- Hex Addr	089E	2206
x"00",	-- Hex Addr	089F	2207
x"00",	-- Hex Addr	08A0	2208
x"00",	-- Hex Addr	08A1	2209
x"00",	-- Hex Addr	08A2	2210
x"00",	-- Hex Addr	08A3	2211
x"00",	-- Hex Addr	08A4	2212
x"00",	-- Hex Addr	08A5	2213
x"00",	-- Hex Addr	08A6	2214
x"00",	-- Hex Addr	08A7	2215
x"00",	-- Hex Addr	08A8	2216
x"00",	-- Hex Addr	08A9	2217
x"00",	-- Hex Addr	08AA	2218
x"00",	-- Hex Addr	08AB	2219
x"00",	-- Hex Addr	08AC	2220
x"00",	-- Hex Addr	08AD	2221
x"00",	-- Hex Addr	08AE	2222
x"00",	-- Hex Addr	08AF	2223
x"00",	-- Hex Addr	08B0	2224
x"00",	-- Hex Addr	08B1	2225
x"00",	-- Hex Addr	08B2	2226
x"00",	-- Hex Addr	08B3	2227
x"00",	-- Hex Addr	08B4	2228
x"00",	-- Hex Addr	08B5	2229
x"00",	-- Hex Addr	08B6	2230
x"00",	-- Hex Addr	08B7	2231
x"00",	-- Hex Addr	08B8	2232
x"00",	-- Hex Addr	08B9	2233
x"00",	-- Hex Addr	08BA	2234
x"00",	-- Hex Addr	08BB	2235
x"00",	-- Hex Addr	08BC	2236
x"00",	-- Hex Addr	08BD	2237
x"00",	-- Hex Addr	08BE	2238
x"00",	-- Hex Addr	08BF	2239
x"00",	-- Hex Addr	08C0	2240
x"00",	-- Hex Addr	08C1	2241
x"00",	-- Hex Addr	08C2	2242
x"00",	-- Hex Addr	08C3	2243
x"00",	-- Hex Addr	08C4	2244
x"00",	-- Hex Addr	08C5	2245
x"00",	-- Hex Addr	08C6	2246
x"00",	-- Hex Addr	08C7	2247
x"00",	-- Hex Addr	08C8	2248
x"00",	-- Hex Addr	08C9	2249
x"00",	-- Hex Addr	08CA	2250
x"00",	-- Hex Addr	08CB	2251
x"00",	-- Hex Addr	08CC	2252
x"00",	-- Hex Addr	08CD	2253
x"00",	-- Hex Addr	08CE	2254
x"00",	-- Hex Addr	08CF	2255
x"00",	-- Hex Addr	08D0	2256
x"00",	-- Hex Addr	08D1	2257
x"00",	-- Hex Addr	08D2	2258
x"00",	-- Hex Addr	08D3	2259
x"00",	-- Hex Addr	08D4	2260
x"00",	-- Hex Addr	08D5	2261
x"00",	-- Hex Addr	08D6	2262
x"00",	-- Hex Addr	08D7	2263
x"00",	-- Hex Addr	08D8	2264
x"00",	-- Hex Addr	08D9	2265
x"00",	-- Hex Addr	08DA	2266
x"00",	-- Hex Addr	08DB	2267
x"00",	-- Hex Addr	08DC	2268
x"00",	-- Hex Addr	08DD	2269
x"00",	-- Hex Addr	08DE	2270
x"00",	-- Hex Addr	08DF	2271
x"00",	-- Hex Addr	08E0	2272
x"00",	-- Hex Addr	08E1	2273
x"00",	-- Hex Addr	08E2	2274
x"00",	-- Hex Addr	08E3	2275
x"00",	-- Hex Addr	08E4	2276
x"00",	-- Hex Addr	08E5	2277
x"00",	-- Hex Addr	08E6	2278
x"00",	-- Hex Addr	08E7	2279
x"00",	-- Hex Addr	08E8	2280
x"00",	-- Hex Addr	08E9	2281
x"00",	-- Hex Addr	08EA	2282
x"00",	-- Hex Addr	08EB	2283
x"00",	-- Hex Addr	08EC	2284
x"00",	-- Hex Addr	08ED	2285
x"00",	-- Hex Addr	08EE	2286
x"00",	-- Hex Addr	08EF	2287
x"00",	-- Hex Addr	08F0	2288
x"00",	-- Hex Addr	08F1	2289
x"00",	-- Hex Addr	08F2	2290
x"00",	-- Hex Addr	08F3	2291
x"00",	-- Hex Addr	08F4	2292
x"00",	-- Hex Addr	08F5	2293
x"00",	-- Hex Addr	08F6	2294
x"00",	-- Hex Addr	08F7	2295
x"00",	-- Hex Addr	08F8	2296
x"00",	-- Hex Addr	08F9	2297
x"00",	-- Hex Addr	08FA	2298
x"00",	-- Hex Addr	08FB	2299
x"00",	-- Hex Addr	08FC	2300
x"00",	-- Hex Addr	08FD	2301
x"00",	-- Hex Addr	08FE	2302
x"00",	-- Hex Addr	08FF	2303
x"00",	-- Hex Addr	0900	2304
x"00",	-- Hex Addr	0901	2305
x"00",	-- Hex Addr	0902	2306
x"00",	-- Hex Addr	0903	2307
x"00",	-- Hex Addr	0904	2308
x"00",	-- Hex Addr	0905	2309
x"00",	-- Hex Addr	0906	2310
x"00",	-- Hex Addr	0907	2311
x"00",	-- Hex Addr	0908	2312
x"00",	-- Hex Addr	0909	2313
x"00",	-- Hex Addr	090A	2314
x"00",	-- Hex Addr	090B	2315
x"00",	-- Hex Addr	090C	2316
x"00",	-- Hex Addr	090D	2317
x"00",	-- Hex Addr	090E	2318
x"00",	-- Hex Addr	090F	2319
x"00",	-- Hex Addr	0910	2320
x"00",	-- Hex Addr	0911	2321
x"00",	-- Hex Addr	0912	2322
x"00",	-- Hex Addr	0913	2323
x"00",	-- Hex Addr	0914	2324
x"00",	-- Hex Addr	0915	2325
x"00",	-- Hex Addr	0916	2326
x"00",	-- Hex Addr	0917	2327
x"00",	-- Hex Addr	0918	2328
x"00",	-- Hex Addr	0919	2329
x"00",	-- Hex Addr	091A	2330
x"00",	-- Hex Addr	091B	2331
x"00",	-- Hex Addr	091C	2332
x"00",	-- Hex Addr	091D	2333
x"00",	-- Hex Addr	091E	2334
x"00",	-- Hex Addr	091F	2335
x"00",	-- Hex Addr	0920	2336
x"00",	-- Hex Addr	0921	2337
x"00",	-- Hex Addr	0922	2338
x"00",	-- Hex Addr	0923	2339
x"00",	-- Hex Addr	0924	2340
x"00",	-- Hex Addr	0925	2341
x"00",	-- Hex Addr	0926	2342
x"00",	-- Hex Addr	0927	2343
x"00",	-- Hex Addr	0928	2344
x"00",	-- Hex Addr	0929	2345
x"00",	-- Hex Addr	092A	2346
x"00",	-- Hex Addr	092B	2347
x"00",	-- Hex Addr	092C	2348
x"00",	-- Hex Addr	092D	2349
x"00",	-- Hex Addr	092E	2350
x"00",	-- Hex Addr	092F	2351
x"00",	-- Hex Addr	0930	2352
x"00",	-- Hex Addr	0931	2353
x"00",	-- Hex Addr	0932	2354
x"00",	-- Hex Addr	0933	2355
x"00",	-- Hex Addr	0934	2356
x"00",	-- Hex Addr	0935	2357
x"00",	-- Hex Addr	0936	2358
x"00",	-- Hex Addr	0937	2359
x"00",	-- Hex Addr	0938	2360
x"00",	-- Hex Addr	0939	2361
x"00",	-- Hex Addr	093A	2362
x"00",	-- Hex Addr	093B	2363
x"00",	-- Hex Addr	093C	2364
x"00",	-- Hex Addr	093D	2365
x"00",	-- Hex Addr	093E	2366
x"00",	-- Hex Addr	093F	2367
x"00",	-- Hex Addr	0940	2368
x"00",	-- Hex Addr	0941	2369
x"00",	-- Hex Addr	0942	2370
x"00",	-- Hex Addr	0943	2371
x"00",	-- Hex Addr	0944	2372
x"00",	-- Hex Addr	0945	2373
x"00",	-- Hex Addr	0946	2374
x"00",	-- Hex Addr	0947	2375
x"00",	-- Hex Addr	0948	2376
x"00",	-- Hex Addr	0949	2377
x"00",	-- Hex Addr	094A	2378
x"00",	-- Hex Addr	094B	2379
x"00",	-- Hex Addr	094C	2380
x"00",	-- Hex Addr	094D	2381
x"00",	-- Hex Addr	094E	2382
x"00",	-- Hex Addr	094F	2383
x"00",	-- Hex Addr	0950	2384
x"00",	-- Hex Addr	0951	2385
x"00",	-- Hex Addr	0952	2386
x"00",	-- Hex Addr	0953	2387
x"00",	-- Hex Addr	0954	2388
x"00",	-- Hex Addr	0955	2389
x"00",	-- Hex Addr	0956	2390
x"00",	-- Hex Addr	0957	2391
x"00",	-- Hex Addr	0958	2392
x"00",	-- Hex Addr	0959	2393
x"00",	-- Hex Addr	095A	2394
x"00",	-- Hex Addr	095B	2395
x"00",	-- Hex Addr	095C	2396
x"00",	-- Hex Addr	095D	2397
x"00",	-- Hex Addr	095E	2398
x"00",	-- Hex Addr	095F	2399
x"00",	-- Hex Addr	0960	2400
x"00",	-- Hex Addr	0961	2401
x"00",	-- Hex Addr	0962	2402
x"00",	-- Hex Addr	0963	2403
x"00",	-- Hex Addr	0964	2404
x"00",	-- Hex Addr	0965	2405
x"00",	-- Hex Addr	0966	2406
x"00",	-- Hex Addr	0967	2407
x"00",	-- Hex Addr	0968	2408
x"00",	-- Hex Addr	0969	2409
x"00",	-- Hex Addr	096A	2410
x"00",	-- Hex Addr	096B	2411
x"00",	-- Hex Addr	096C	2412
x"00",	-- Hex Addr	096D	2413
x"00",	-- Hex Addr	096E	2414
x"00",	-- Hex Addr	096F	2415
x"00",	-- Hex Addr	0970	2416
x"00",	-- Hex Addr	0971	2417
x"00",	-- Hex Addr	0972	2418
x"00",	-- Hex Addr	0973	2419
x"00",	-- Hex Addr	0974	2420
x"00",	-- Hex Addr	0975	2421
x"00",	-- Hex Addr	0976	2422
x"00",	-- Hex Addr	0977	2423
x"00",	-- Hex Addr	0978	2424
x"00",	-- Hex Addr	0979	2425
x"00",	-- Hex Addr	097A	2426
x"00",	-- Hex Addr	097B	2427
x"00",	-- Hex Addr	097C	2428
x"00",	-- Hex Addr	097D	2429
x"00",	-- Hex Addr	097E	2430
x"00",	-- Hex Addr	097F	2431
x"00",	-- Hex Addr	0980	2432
x"00",	-- Hex Addr	0981	2433
x"00",	-- Hex Addr	0982	2434
x"00",	-- Hex Addr	0983	2435
x"00",	-- Hex Addr	0984	2436
x"00",	-- Hex Addr	0985	2437
x"00",	-- Hex Addr	0986	2438
x"00",	-- Hex Addr	0987	2439
x"00",	-- Hex Addr	0988	2440
x"00",	-- Hex Addr	0989	2441
x"00",	-- Hex Addr	098A	2442
x"00",	-- Hex Addr	098B	2443
x"00",	-- Hex Addr	098C	2444
x"00",	-- Hex Addr	098D	2445
x"00",	-- Hex Addr	098E	2446
x"00",	-- Hex Addr	098F	2447
x"00",	-- Hex Addr	0990	2448
x"00",	-- Hex Addr	0991	2449
x"00",	-- Hex Addr	0992	2450
x"00",	-- Hex Addr	0993	2451
x"00",	-- Hex Addr	0994	2452
x"00",	-- Hex Addr	0995	2453
x"00",	-- Hex Addr	0996	2454
x"00",	-- Hex Addr	0997	2455
x"00",	-- Hex Addr	0998	2456
x"00",	-- Hex Addr	0999	2457
x"00",	-- Hex Addr	099A	2458
x"00",	-- Hex Addr	099B	2459
x"00",	-- Hex Addr	099C	2460
x"00",	-- Hex Addr	099D	2461
x"00",	-- Hex Addr	099E	2462
x"00",	-- Hex Addr	099F	2463
x"00",	-- Hex Addr	09A0	2464
x"00",	-- Hex Addr	09A1	2465
x"00",	-- Hex Addr	09A2	2466
x"00",	-- Hex Addr	09A3	2467
x"00",	-- Hex Addr	09A4	2468
x"00",	-- Hex Addr	09A5	2469
x"00",	-- Hex Addr	09A6	2470
x"00",	-- Hex Addr	09A7	2471
x"00",	-- Hex Addr	09A8	2472
x"00",	-- Hex Addr	09A9	2473
x"00",	-- Hex Addr	09AA	2474
x"00",	-- Hex Addr	09AB	2475
x"00",	-- Hex Addr	09AC	2476
x"00",	-- Hex Addr	09AD	2477
x"00",	-- Hex Addr	09AE	2478
x"00",	-- Hex Addr	09AF	2479
x"00",	-- Hex Addr	09B0	2480
x"00",	-- Hex Addr	09B1	2481
x"00",	-- Hex Addr	09B2	2482
x"00",	-- Hex Addr	09B3	2483
x"00",	-- Hex Addr	09B4	2484
x"00",	-- Hex Addr	09B5	2485
x"00",	-- Hex Addr	09B6	2486
x"00",	-- Hex Addr	09B7	2487
x"00",	-- Hex Addr	09B8	2488
x"00",	-- Hex Addr	09B9	2489
x"00",	-- Hex Addr	09BA	2490
x"00",	-- Hex Addr	09BB	2491
x"00",	-- Hex Addr	09BC	2492
x"00",	-- Hex Addr	09BD	2493
x"00",	-- Hex Addr	09BE	2494
x"00",	-- Hex Addr	09BF	2495
x"00",	-- Hex Addr	09C0	2496
x"00",	-- Hex Addr	09C1	2497
x"00",	-- Hex Addr	09C2	2498
x"00",	-- Hex Addr	09C3	2499
x"00",	-- Hex Addr	09C4	2500
x"00",	-- Hex Addr	09C5	2501
x"00",	-- Hex Addr	09C6	2502
x"00",	-- Hex Addr	09C7	2503
x"00",	-- Hex Addr	09C8	2504
x"00",	-- Hex Addr	09C9	2505
x"00",	-- Hex Addr	09CA	2506
x"00",	-- Hex Addr	09CB	2507
x"00",	-- Hex Addr	09CC	2508
x"00",	-- Hex Addr	09CD	2509
x"00",	-- Hex Addr	09CE	2510
x"00",	-- Hex Addr	09CF	2511
x"00",	-- Hex Addr	09D0	2512
x"00",	-- Hex Addr	09D1	2513
x"00",	-- Hex Addr	09D2	2514
x"00",	-- Hex Addr	09D3	2515
x"00",	-- Hex Addr	09D4	2516
x"00",	-- Hex Addr	09D5	2517
x"00",	-- Hex Addr	09D6	2518
x"00",	-- Hex Addr	09D7	2519
x"00",	-- Hex Addr	09D8	2520
x"00",	-- Hex Addr	09D9	2521
x"00",	-- Hex Addr	09DA	2522
x"00",	-- Hex Addr	09DB	2523
x"00",	-- Hex Addr	09DC	2524
x"00",	-- Hex Addr	09DD	2525
x"00",	-- Hex Addr	09DE	2526
x"00",	-- Hex Addr	09DF	2527
x"00",	-- Hex Addr	09E0	2528
x"00",	-- Hex Addr	09E1	2529
x"00",	-- Hex Addr	09E2	2530
x"00",	-- Hex Addr	09E3	2531
x"00",	-- Hex Addr	09E4	2532
x"00",	-- Hex Addr	09E5	2533
x"00",	-- Hex Addr	09E6	2534
x"00",	-- Hex Addr	09E7	2535
x"00",	-- Hex Addr	09E8	2536
x"00",	-- Hex Addr	09E9	2537
x"00",	-- Hex Addr	09EA	2538
x"00",	-- Hex Addr	09EB	2539
x"00",	-- Hex Addr	09EC	2540
x"00",	-- Hex Addr	09ED	2541
x"00",	-- Hex Addr	09EE	2542
x"00",	-- Hex Addr	09EF	2543
x"00",	-- Hex Addr	09F0	2544
x"00",	-- Hex Addr	09F1	2545
x"00",	-- Hex Addr	09F2	2546
x"00",	-- Hex Addr	09F3	2547
x"00",	-- Hex Addr	09F4	2548
x"00",	-- Hex Addr	09F5	2549
x"00",	-- Hex Addr	09F6	2550
x"00",	-- Hex Addr	09F7	2551
x"00",	-- Hex Addr	09F8	2552
x"00",	-- Hex Addr	09F9	2553
x"00",	-- Hex Addr	09FA	2554
x"00",	-- Hex Addr	09FB	2555
x"00",	-- Hex Addr	09FC	2556
x"00",	-- Hex Addr	09FD	2557
x"00",	-- Hex Addr	09FE	2558
x"00",	-- Hex Addr	09FF	2559
x"00",	-- Hex Addr	0A00	2560
x"00",	-- Hex Addr	0A01	2561
x"00",	-- Hex Addr	0A02	2562
x"00",	-- Hex Addr	0A03	2563
x"00",	-- Hex Addr	0A04	2564
x"00",	-- Hex Addr	0A05	2565
x"00",	-- Hex Addr	0A06	2566
x"00",	-- Hex Addr	0A07	2567
x"00",	-- Hex Addr	0A08	2568
x"00",	-- Hex Addr	0A09	2569
x"00",	-- Hex Addr	0A0A	2570
x"00",	-- Hex Addr	0A0B	2571
x"00",	-- Hex Addr	0A0C	2572
x"00",	-- Hex Addr	0A0D	2573
x"00",	-- Hex Addr	0A0E	2574
x"00",	-- Hex Addr	0A0F	2575
x"00",	-- Hex Addr	0A10	2576
x"00",	-- Hex Addr	0A11	2577
x"00",	-- Hex Addr	0A12	2578
x"00",	-- Hex Addr	0A13	2579
x"00",	-- Hex Addr	0A14	2580
x"00",	-- Hex Addr	0A15	2581
x"00",	-- Hex Addr	0A16	2582
x"00",	-- Hex Addr	0A17	2583
x"00",	-- Hex Addr	0A18	2584
x"00",	-- Hex Addr	0A19	2585
x"00",	-- Hex Addr	0A1A	2586
x"00",	-- Hex Addr	0A1B	2587
x"00",	-- Hex Addr	0A1C	2588
x"00",	-- Hex Addr	0A1D	2589
x"00",	-- Hex Addr	0A1E	2590
x"00",	-- Hex Addr	0A1F	2591
x"00",	-- Hex Addr	0A20	2592
x"00",	-- Hex Addr	0A21	2593
x"00",	-- Hex Addr	0A22	2594
x"00",	-- Hex Addr	0A23	2595
x"00",	-- Hex Addr	0A24	2596
x"00",	-- Hex Addr	0A25	2597
x"00",	-- Hex Addr	0A26	2598
x"00",	-- Hex Addr	0A27	2599
x"00",	-- Hex Addr	0A28	2600
x"00",	-- Hex Addr	0A29	2601
x"00",	-- Hex Addr	0A2A	2602
x"00",	-- Hex Addr	0A2B	2603
x"00",	-- Hex Addr	0A2C	2604
x"00",	-- Hex Addr	0A2D	2605
x"00",	-- Hex Addr	0A2E	2606
x"00",	-- Hex Addr	0A2F	2607
x"00",	-- Hex Addr	0A30	2608
x"00",	-- Hex Addr	0A31	2609
x"00",	-- Hex Addr	0A32	2610
x"00",	-- Hex Addr	0A33	2611
x"00",	-- Hex Addr	0A34	2612
x"00",	-- Hex Addr	0A35	2613
x"00",	-- Hex Addr	0A36	2614
x"00",	-- Hex Addr	0A37	2615
x"00",	-- Hex Addr	0A38	2616
x"00",	-- Hex Addr	0A39	2617
x"00",	-- Hex Addr	0A3A	2618
x"00",	-- Hex Addr	0A3B	2619
x"00",	-- Hex Addr	0A3C	2620
x"00",	-- Hex Addr	0A3D	2621
x"00",	-- Hex Addr	0A3E	2622
x"00",	-- Hex Addr	0A3F	2623
x"00",	-- Hex Addr	0A40	2624
x"00",	-- Hex Addr	0A41	2625
x"00",	-- Hex Addr	0A42	2626
x"00",	-- Hex Addr	0A43	2627
x"00",	-- Hex Addr	0A44	2628
x"00",	-- Hex Addr	0A45	2629
x"00",	-- Hex Addr	0A46	2630
x"00",	-- Hex Addr	0A47	2631
x"00",	-- Hex Addr	0A48	2632
x"00",	-- Hex Addr	0A49	2633
x"00",	-- Hex Addr	0A4A	2634
x"00",	-- Hex Addr	0A4B	2635
x"00",	-- Hex Addr	0A4C	2636
x"00",	-- Hex Addr	0A4D	2637
x"00",	-- Hex Addr	0A4E	2638
x"00",	-- Hex Addr	0A4F	2639
x"00",	-- Hex Addr	0A50	2640
x"00",	-- Hex Addr	0A51	2641
x"00",	-- Hex Addr	0A52	2642
x"00",	-- Hex Addr	0A53	2643
x"00",	-- Hex Addr	0A54	2644
x"00",	-- Hex Addr	0A55	2645
x"00",	-- Hex Addr	0A56	2646
x"00",	-- Hex Addr	0A57	2647
x"00",	-- Hex Addr	0A58	2648
x"00",	-- Hex Addr	0A59	2649
x"00",	-- Hex Addr	0A5A	2650
x"00",	-- Hex Addr	0A5B	2651
x"00",	-- Hex Addr	0A5C	2652
x"00",	-- Hex Addr	0A5D	2653
x"00",	-- Hex Addr	0A5E	2654
x"00",	-- Hex Addr	0A5F	2655
x"00",	-- Hex Addr	0A60	2656
x"00",	-- Hex Addr	0A61	2657
x"00",	-- Hex Addr	0A62	2658
x"00",	-- Hex Addr	0A63	2659
x"00",	-- Hex Addr	0A64	2660
x"00",	-- Hex Addr	0A65	2661
x"00",	-- Hex Addr	0A66	2662
x"00",	-- Hex Addr	0A67	2663
x"00",	-- Hex Addr	0A68	2664
x"00",	-- Hex Addr	0A69	2665
x"00",	-- Hex Addr	0A6A	2666
x"00",	-- Hex Addr	0A6B	2667
x"00",	-- Hex Addr	0A6C	2668
x"00",	-- Hex Addr	0A6D	2669
x"00",	-- Hex Addr	0A6E	2670
x"00",	-- Hex Addr	0A6F	2671
x"00",	-- Hex Addr	0A70	2672
x"00",	-- Hex Addr	0A71	2673
x"00",	-- Hex Addr	0A72	2674
x"00",	-- Hex Addr	0A73	2675
x"00",	-- Hex Addr	0A74	2676
x"00",	-- Hex Addr	0A75	2677
x"00",	-- Hex Addr	0A76	2678
x"00",	-- Hex Addr	0A77	2679
x"00",	-- Hex Addr	0A78	2680
x"00",	-- Hex Addr	0A79	2681
x"00",	-- Hex Addr	0A7A	2682
x"00",	-- Hex Addr	0A7B	2683
x"00",	-- Hex Addr	0A7C	2684
x"00",	-- Hex Addr	0A7D	2685
x"00",	-- Hex Addr	0A7E	2686
x"00",	-- Hex Addr	0A7F	2687
x"00",	-- Hex Addr	0A80	2688
x"00",	-- Hex Addr	0A81	2689
x"00",	-- Hex Addr	0A82	2690
x"00",	-- Hex Addr	0A83	2691
x"00",	-- Hex Addr	0A84	2692
x"00",	-- Hex Addr	0A85	2693
x"00",	-- Hex Addr	0A86	2694
x"00",	-- Hex Addr	0A87	2695
x"00",	-- Hex Addr	0A88	2696
x"00",	-- Hex Addr	0A89	2697
x"00",	-- Hex Addr	0A8A	2698
x"00",	-- Hex Addr	0A8B	2699
x"00",	-- Hex Addr	0A8C	2700
x"00",	-- Hex Addr	0A8D	2701
x"00",	-- Hex Addr	0A8E	2702
x"00",	-- Hex Addr	0A8F	2703
x"00",	-- Hex Addr	0A90	2704
x"00",	-- Hex Addr	0A91	2705
x"00",	-- Hex Addr	0A92	2706
x"00",	-- Hex Addr	0A93	2707
x"00",	-- Hex Addr	0A94	2708
x"00",	-- Hex Addr	0A95	2709
x"00",	-- Hex Addr	0A96	2710
x"00",	-- Hex Addr	0A97	2711
x"00",	-- Hex Addr	0A98	2712
x"00",	-- Hex Addr	0A99	2713
x"00",	-- Hex Addr	0A9A	2714
x"00",	-- Hex Addr	0A9B	2715
x"00",	-- Hex Addr	0A9C	2716
x"00",	-- Hex Addr	0A9D	2717
x"00",	-- Hex Addr	0A9E	2718
x"00",	-- Hex Addr	0A9F	2719
x"00",	-- Hex Addr	0AA0	2720
x"00",	-- Hex Addr	0AA1	2721
x"00",	-- Hex Addr	0AA2	2722
x"00",	-- Hex Addr	0AA3	2723
x"00",	-- Hex Addr	0AA4	2724
x"00",	-- Hex Addr	0AA5	2725
x"00",	-- Hex Addr	0AA6	2726
x"00",	-- Hex Addr	0AA7	2727
x"00",	-- Hex Addr	0AA8	2728
x"00",	-- Hex Addr	0AA9	2729
x"00",	-- Hex Addr	0AAA	2730
x"00",	-- Hex Addr	0AAB	2731
x"00",	-- Hex Addr	0AAC	2732
x"00",	-- Hex Addr	0AAD	2733
x"00",	-- Hex Addr	0AAE	2734
x"00",	-- Hex Addr	0AAF	2735
x"00",	-- Hex Addr	0AB0	2736
x"00",	-- Hex Addr	0AB1	2737
x"00",	-- Hex Addr	0AB2	2738
x"00",	-- Hex Addr	0AB3	2739
x"00",	-- Hex Addr	0AB4	2740
x"00",	-- Hex Addr	0AB5	2741
x"00",	-- Hex Addr	0AB6	2742
x"00",	-- Hex Addr	0AB7	2743
x"00",	-- Hex Addr	0AB8	2744
x"00",	-- Hex Addr	0AB9	2745
x"00",	-- Hex Addr	0ABA	2746
x"00",	-- Hex Addr	0ABB	2747
x"00",	-- Hex Addr	0ABC	2748
x"00",	-- Hex Addr	0ABD	2749
x"00",	-- Hex Addr	0ABE	2750
x"00",	-- Hex Addr	0ABF	2751
x"00",	-- Hex Addr	0AC0	2752
x"00",	-- Hex Addr	0AC1	2753
x"00",	-- Hex Addr	0AC2	2754
x"00",	-- Hex Addr	0AC3	2755
x"00",	-- Hex Addr	0AC4	2756
x"00",	-- Hex Addr	0AC5	2757
x"00",	-- Hex Addr	0AC6	2758
x"00",	-- Hex Addr	0AC7	2759
x"00",	-- Hex Addr	0AC8	2760
x"00",	-- Hex Addr	0AC9	2761
x"00",	-- Hex Addr	0ACA	2762
x"00",	-- Hex Addr	0ACB	2763
x"00",	-- Hex Addr	0ACC	2764
x"00",	-- Hex Addr	0ACD	2765
x"00",	-- Hex Addr	0ACE	2766
x"00",	-- Hex Addr	0ACF	2767
x"00",	-- Hex Addr	0AD0	2768
x"00",	-- Hex Addr	0AD1	2769
x"00",	-- Hex Addr	0AD2	2770
x"00",	-- Hex Addr	0AD3	2771
x"00",	-- Hex Addr	0AD4	2772
x"00",	-- Hex Addr	0AD5	2773
x"00",	-- Hex Addr	0AD6	2774
x"00",	-- Hex Addr	0AD7	2775
x"00",	-- Hex Addr	0AD8	2776
x"00",	-- Hex Addr	0AD9	2777
x"00",	-- Hex Addr	0ADA	2778
x"00",	-- Hex Addr	0ADB	2779
x"00",	-- Hex Addr	0ADC	2780
x"00",	-- Hex Addr	0ADD	2781
x"00",	-- Hex Addr	0ADE	2782
x"00",	-- Hex Addr	0ADF	2783
x"00",	-- Hex Addr	0AE0	2784
x"00",	-- Hex Addr	0AE1	2785
x"00",	-- Hex Addr	0AE2	2786
x"00",	-- Hex Addr	0AE3	2787
x"00",	-- Hex Addr	0AE4	2788
x"00",	-- Hex Addr	0AE5	2789
x"00",	-- Hex Addr	0AE6	2790
x"00",	-- Hex Addr	0AE7	2791
x"00",	-- Hex Addr	0AE8	2792
x"00",	-- Hex Addr	0AE9	2793
x"00",	-- Hex Addr	0AEA	2794
x"00",	-- Hex Addr	0AEB	2795
x"00",	-- Hex Addr	0AEC	2796
x"00",	-- Hex Addr	0AED	2797
x"00",	-- Hex Addr	0AEE	2798
x"00",	-- Hex Addr	0AEF	2799
x"00",	-- Hex Addr	0AF0	2800
x"00",	-- Hex Addr	0AF1	2801
x"00",	-- Hex Addr	0AF2	2802
x"00",	-- Hex Addr	0AF3	2803
x"00",	-- Hex Addr	0AF4	2804
x"00",	-- Hex Addr	0AF5	2805
x"00",	-- Hex Addr	0AF6	2806
x"00",	-- Hex Addr	0AF7	2807
x"00",	-- Hex Addr	0AF8	2808
x"00",	-- Hex Addr	0AF9	2809
x"00",	-- Hex Addr	0AFA	2810
x"00",	-- Hex Addr	0AFB	2811
x"00",	-- Hex Addr	0AFC	2812
x"00",	-- Hex Addr	0AFD	2813
x"00",	-- Hex Addr	0AFE	2814
x"00",	-- Hex Addr	0AFF	2815
x"00",	-- Hex Addr	0B00	2816
x"00",	-- Hex Addr	0B01	2817
x"00",	-- Hex Addr	0B02	2818
x"00",	-- Hex Addr	0B03	2819
x"00",	-- Hex Addr	0B04	2820
x"00",	-- Hex Addr	0B05	2821
x"00",	-- Hex Addr	0B06	2822
x"00",	-- Hex Addr	0B07	2823
x"00",	-- Hex Addr	0B08	2824
x"00",	-- Hex Addr	0B09	2825
x"00",	-- Hex Addr	0B0A	2826
x"00",	-- Hex Addr	0B0B	2827
x"00",	-- Hex Addr	0B0C	2828
x"00",	-- Hex Addr	0B0D	2829
x"00",	-- Hex Addr	0B0E	2830
x"00",	-- Hex Addr	0B0F	2831
x"00",	-- Hex Addr	0B10	2832
x"00",	-- Hex Addr	0B11	2833
x"00",	-- Hex Addr	0B12	2834
x"00",	-- Hex Addr	0B13	2835
x"00",	-- Hex Addr	0B14	2836
x"00",	-- Hex Addr	0B15	2837
x"00",	-- Hex Addr	0B16	2838
x"00",	-- Hex Addr	0B17	2839
x"00",	-- Hex Addr	0B18	2840
x"00",	-- Hex Addr	0B19	2841
x"00",	-- Hex Addr	0B1A	2842
x"00",	-- Hex Addr	0B1B	2843
x"00",	-- Hex Addr	0B1C	2844
x"00",	-- Hex Addr	0B1D	2845
x"00",	-- Hex Addr	0B1E	2846
x"00",	-- Hex Addr	0B1F	2847
x"00",	-- Hex Addr	0B20	2848
x"00",	-- Hex Addr	0B21	2849
x"00",	-- Hex Addr	0B22	2850
x"00",	-- Hex Addr	0B23	2851
x"00",	-- Hex Addr	0B24	2852
x"00",	-- Hex Addr	0B25	2853
x"00",	-- Hex Addr	0B26	2854
x"00",	-- Hex Addr	0B27	2855
x"00",	-- Hex Addr	0B28	2856
x"00",	-- Hex Addr	0B29	2857
x"00",	-- Hex Addr	0B2A	2858
x"00",	-- Hex Addr	0B2B	2859
x"00",	-- Hex Addr	0B2C	2860
x"00",	-- Hex Addr	0B2D	2861
x"00",	-- Hex Addr	0B2E	2862
x"00",	-- Hex Addr	0B2F	2863
x"00",	-- Hex Addr	0B30	2864
x"00",	-- Hex Addr	0B31	2865
x"00",	-- Hex Addr	0B32	2866
x"00",	-- Hex Addr	0B33	2867
x"00",	-- Hex Addr	0B34	2868
x"00",	-- Hex Addr	0B35	2869
x"00",	-- Hex Addr	0B36	2870
x"00",	-- Hex Addr	0B37	2871
x"00",	-- Hex Addr	0B38	2872
x"00",	-- Hex Addr	0B39	2873
x"00",	-- Hex Addr	0B3A	2874
x"00",	-- Hex Addr	0B3B	2875
x"00",	-- Hex Addr	0B3C	2876
x"00",	-- Hex Addr	0B3D	2877
x"00",	-- Hex Addr	0B3E	2878
x"00",	-- Hex Addr	0B3F	2879
x"00",	-- Hex Addr	0B40	2880
x"00",	-- Hex Addr	0B41	2881
x"00",	-- Hex Addr	0B42	2882
x"00",	-- Hex Addr	0B43	2883
x"00",	-- Hex Addr	0B44	2884
x"00",	-- Hex Addr	0B45	2885
x"00",	-- Hex Addr	0B46	2886
x"00",	-- Hex Addr	0B47	2887
x"00",	-- Hex Addr	0B48	2888
x"00",	-- Hex Addr	0B49	2889
x"00",	-- Hex Addr	0B4A	2890
x"00",	-- Hex Addr	0B4B	2891
x"00",	-- Hex Addr	0B4C	2892
x"00",	-- Hex Addr	0B4D	2893
x"00",	-- Hex Addr	0B4E	2894
x"00",	-- Hex Addr	0B4F	2895
x"00",	-- Hex Addr	0B50	2896
x"00",	-- Hex Addr	0B51	2897
x"00",	-- Hex Addr	0B52	2898
x"00",	-- Hex Addr	0B53	2899
x"00",	-- Hex Addr	0B54	2900
x"00",	-- Hex Addr	0B55	2901
x"00",	-- Hex Addr	0B56	2902
x"00",	-- Hex Addr	0B57	2903
x"00",	-- Hex Addr	0B58	2904
x"00",	-- Hex Addr	0B59	2905
x"00",	-- Hex Addr	0B5A	2906
x"00",	-- Hex Addr	0B5B	2907
x"00",	-- Hex Addr	0B5C	2908
x"00",	-- Hex Addr	0B5D	2909
x"00",	-- Hex Addr	0B5E	2910
x"00",	-- Hex Addr	0B5F	2911
x"00",	-- Hex Addr	0B60	2912
x"00",	-- Hex Addr	0B61	2913
x"00",	-- Hex Addr	0B62	2914
x"00",	-- Hex Addr	0B63	2915
x"00",	-- Hex Addr	0B64	2916
x"00",	-- Hex Addr	0B65	2917
x"00",	-- Hex Addr	0B66	2918
x"00",	-- Hex Addr	0B67	2919
x"00",	-- Hex Addr	0B68	2920
x"00",	-- Hex Addr	0B69	2921
x"00",	-- Hex Addr	0B6A	2922
x"00",	-- Hex Addr	0B6B	2923
x"00",	-- Hex Addr	0B6C	2924
x"00",	-- Hex Addr	0B6D	2925
x"00",	-- Hex Addr	0B6E	2926
x"00",	-- Hex Addr	0B6F	2927
x"00",	-- Hex Addr	0B70	2928
x"00",	-- Hex Addr	0B71	2929
x"00",	-- Hex Addr	0B72	2930
x"00",	-- Hex Addr	0B73	2931
x"00",	-- Hex Addr	0B74	2932
x"00",	-- Hex Addr	0B75	2933
x"00",	-- Hex Addr	0B76	2934
x"00",	-- Hex Addr	0B77	2935
x"00",	-- Hex Addr	0B78	2936
x"00",	-- Hex Addr	0B79	2937
x"00",	-- Hex Addr	0B7A	2938
x"00",	-- Hex Addr	0B7B	2939
x"00",	-- Hex Addr	0B7C	2940
x"00",	-- Hex Addr	0B7D	2941
x"00",	-- Hex Addr	0B7E	2942
x"00",	-- Hex Addr	0B7F	2943
x"00",	-- Hex Addr	0B80	2944
x"00",	-- Hex Addr	0B81	2945
x"00",	-- Hex Addr	0B82	2946
x"00",	-- Hex Addr	0B83	2947
x"00",	-- Hex Addr	0B84	2948
x"00",	-- Hex Addr	0B85	2949
x"00",	-- Hex Addr	0B86	2950
x"00",	-- Hex Addr	0B87	2951
x"00",	-- Hex Addr	0B88	2952
x"00",	-- Hex Addr	0B89	2953
x"00",	-- Hex Addr	0B8A	2954
x"00",	-- Hex Addr	0B8B	2955
x"00",	-- Hex Addr	0B8C	2956
x"00",	-- Hex Addr	0B8D	2957
x"00",	-- Hex Addr	0B8E	2958
x"00",	-- Hex Addr	0B8F	2959
x"00",	-- Hex Addr	0B90	2960
x"00",	-- Hex Addr	0B91	2961
x"00",	-- Hex Addr	0B92	2962
x"00",	-- Hex Addr	0B93	2963
x"00",	-- Hex Addr	0B94	2964
x"00",	-- Hex Addr	0B95	2965
x"00",	-- Hex Addr	0B96	2966
x"00",	-- Hex Addr	0B97	2967
x"00",	-- Hex Addr	0B98	2968
x"00",	-- Hex Addr	0B99	2969
x"00",	-- Hex Addr	0B9A	2970
x"00",	-- Hex Addr	0B9B	2971
x"00",	-- Hex Addr	0B9C	2972
x"00",	-- Hex Addr	0B9D	2973
x"00",	-- Hex Addr	0B9E	2974
x"00",	-- Hex Addr	0B9F	2975
x"00",	-- Hex Addr	0BA0	2976
x"00",	-- Hex Addr	0BA1	2977
x"00",	-- Hex Addr	0BA2	2978
x"00",	-- Hex Addr	0BA3	2979
x"00",	-- Hex Addr	0BA4	2980
x"00",	-- Hex Addr	0BA5	2981
x"00",	-- Hex Addr	0BA6	2982
x"00",	-- Hex Addr	0BA7	2983
x"00",	-- Hex Addr	0BA8	2984
x"00",	-- Hex Addr	0BA9	2985
x"00",	-- Hex Addr	0BAA	2986
x"00",	-- Hex Addr	0BAB	2987
x"00",	-- Hex Addr	0BAC	2988
x"00",	-- Hex Addr	0BAD	2989
x"00",	-- Hex Addr	0BAE	2990
x"00",	-- Hex Addr	0BAF	2991
x"00",	-- Hex Addr	0BB0	2992
x"00",	-- Hex Addr	0BB1	2993
x"00",	-- Hex Addr	0BB2	2994
x"00",	-- Hex Addr	0BB3	2995
x"00",	-- Hex Addr	0BB4	2996
x"00",	-- Hex Addr	0BB5	2997
x"00",	-- Hex Addr	0BB6	2998
x"00",	-- Hex Addr	0BB7	2999
x"00",	-- Hex Addr	0BB8	3000
x"00",	-- Hex Addr	0BB9	3001
x"00",	-- Hex Addr	0BBA	3002
x"00",	-- Hex Addr	0BBB	3003
x"00",	-- Hex Addr	0BBC	3004
x"00",	-- Hex Addr	0BBD	3005
x"00",	-- Hex Addr	0BBE	3006
x"00",	-- Hex Addr	0BBF	3007
x"00",	-- Hex Addr	0BC0	3008
x"00",	-- Hex Addr	0BC1	3009
x"00",	-- Hex Addr	0BC2	3010
x"00",	-- Hex Addr	0BC3	3011
x"00",	-- Hex Addr	0BC4	3012
x"00",	-- Hex Addr	0BC5	3013
x"00",	-- Hex Addr	0BC6	3014
x"00",	-- Hex Addr	0BC7	3015
x"00",	-- Hex Addr	0BC8	3016
x"00",	-- Hex Addr	0BC9	3017
x"00",	-- Hex Addr	0BCA	3018
x"00",	-- Hex Addr	0BCB	3019
x"00",	-- Hex Addr	0BCC	3020
x"00",	-- Hex Addr	0BCD	3021
x"00",	-- Hex Addr	0BCE	3022
x"00",	-- Hex Addr	0BCF	3023
x"00",	-- Hex Addr	0BD0	3024
x"00",	-- Hex Addr	0BD1	3025
x"00",	-- Hex Addr	0BD2	3026
x"00",	-- Hex Addr	0BD3	3027
x"00",	-- Hex Addr	0BD4	3028
x"00",	-- Hex Addr	0BD5	3029
x"00",	-- Hex Addr	0BD6	3030
x"00",	-- Hex Addr	0BD7	3031
x"00",	-- Hex Addr	0BD8	3032
x"00",	-- Hex Addr	0BD9	3033
x"00",	-- Hex Addr	0BDA	3034
x"00",	-- Hex Addr	0BDB	3035
x"00",	-- Hex Addr	0BDC	3036
x"00",	-- Hex Addr	0BDD	3037
x"00",	-- Hex Addr	0BDE	3038
x"00",	-- Hex Addr	0BDF	3039
x"00",	-- Hex Addr	0BE0	3040
x"00",	-- Hex Addr	0BE1	3041
x"00",	-- Hex Addr	0BE2	3042
x"00",	-- Hex Addr	0BE3	3043
x"00",	-- Hex Addr	0BE4	3044
x"00",	-- Hex Addr	0BE5	3045
x"00",	-- Hex Addr	0BE6	3046
x"00",	-- Hex Addr	0BE7	3047
x"00",	-- Hex Addr	0BE8	3048
x"00",	-- Hex Addr	0BE9	3049
x"00",	-- Hex Addr	0BEA	3050
x"00",	-- Hex Addr	0BEB	3051
x"00",	-- Hex Addr	0BEC	3052
x"00",	-- Hex Addr	0BED	3053
x"00",	-- Hex Addr	0BEE	3054
x"00",	-- Hex Addr	0BEF	3055
x"00",	-- Hex Addr	0BF0	3056
x"00",	-- Hex Addr	0BF1	3057
x"00",	-- Hex Addr	0BF2	3058
x"00",	-- Hex Addr	0BF3	3059
x"00",	-- Hex Addr	0BF4	3060
x"00",	-- Hex Addr	0BF5	3061
x"00",	-- Hex Addr	0BF6	3062
x"00",	-- Hex Addr	0BF7	3063
x"00",	-- Hex Addr	0BF8	3064
x"00",	-- Hex Addr	0BF9	3065
x"00",	-- Hex Addr	0BFA	3066
x"00",	-- Hex Addr	0BFB	3067
x"00",	-- Hex Addr	0BFC	3068
x"00",	-- Hex Addr	0BFD	3069
x"00",	-- Hex Addr	0BFE	3070
x"00",	-- Hex Addr	0BFF	3071
x"00",	-- Hex Addr	0C00	3072
x"00",	-- Hex Addr	0C01	3073
x"00",	-- Hex Addr	0C02	3074
x"00",	-- Hex Addr	0C03	3075
x"00",	-- Hex Addr	0C04	3076
x"00",	-- Hex Addr	0C05	3077
x"00",	-- Hex Addr	0C06	3078
x"00",	-- Hex Addr	0C07	3079
x"00",	-- Hex Addr	0C08	3080
x"00",	-- Hex Addr	0C09	3081
x"00",	-- Hex Addr	0C0A	3082
x"00",	-- Hex Addr	0C0B	3083
x"00",	-- Hex Addr	0C0C	3084
x"00",	-- Hex Addr	0C0D	3085
x"00",	-- Hex Addr	0C0E	3086
x"00",	-- Hex Addr	0C0F	3087
x"00",	-- Hex Addr	0C10	3088
x"00",	-- Hex Addr	0C11	3089
x"00",	-- Hex Addr	0C12	3090
x"00",	-- Hex Addr	0C13	3091
x"00",	-- Hex Addr	0C14	3092
x"00",	-- Hex Addr	0C15	3093
x"00",	-- Hex Addr	0C16	3094
x"00",	-- Hex Addr	0C17	3095
x"00",	-- Hex Addr	0C18	3096
x"00",	-- Hex Addr	0C19	3097
x"00",	-- Hex Addr	0C1A	3098
x"00",	-- Hex Addr	0C1B	3099
x"00",	-- Hex Addr	0C1C	3100
x"00",	-- Hex Addr	0C1D	3101
x"00",	-- Hex Addr	0C1E	3102
x"00",	-- Hex Addr	0C1F	3103
x"00",	-- Hex Addr	0C20	3104
x"00",	-- Hex Addr	0C21	3105
x"00",	-- Hex Addr	0C22	3106
x"00",	-- Hex Addr	0C23	3107
x"00",	-- Hex Addr	0C24	3108
x"00",	-- Hex Addr	0C25	3109
x"00",	-- Hex Addr	0C26	3110
x"00",	-- Hex Addr	0C27	3111
x"00",	-- Hex Addr	0C28	3112
x"00",	-- Hex Addr	0C29	3113
x"00",	-- Hex Addr	0C2A	3114
x"00",	-- Hex Addr	0C2B	3115
x"00",	-- Hex Addr	0C2C	3116
x"00",	-- Hex Addr	0C2D	3117
x"00",	-- Hex Addr	0C2E	3118
x"00",	-- Hex Addr	0C2F	3119
x"00",	-- Hex Addr	0C30	3120
x"00",	-- Hex Addr	0C31	3121
x"00",	-- Hex Addr	0C32	3122
x"00",	-- Hex Addr	0C33	3123
x"00",	-- Hex Addr	0C34	3124
x"00",	-- Hex Addr	0C35	3125
x"00",	-- Hex Addr	0C36	3126
x"00",	-- Hex Addr	0C37	3127
x"00",	-- Hex Addr	0C38	3128
x"00",	-- Hex Addr	0C39	3129
x"00",	-- Hex Addr	0C3A	3130
x"00",	-- Hex Addr	0C3B	3131
x"00",	-- Hex Addr	0C3C	3132
x"00",	-- Hex Addr	0C3D	3133
x"00",	-- Hex Addr	0C3E	3134
x"00",	-- Hex Addr	0C3F	3135
x"00",	-- Hex Addr	0C40	3136
x"00",	-- Hex Addr	0C41	3137
x"00",	-- Hex Addr	0C42	3138
x"00",	-- Hex Addr	0C43	3139
x"00",	-- Hex Addr	0C44	3140
x"00",	-- Hex Addr	0C45	3141
x"00",	-- Hex Addr	0C46	3142
x"00",	-- Hex Addr	0C47	3143
x"00",	-- Hex Addr	0C48	3144
x"00",	-- Hex Addr	0C49	3145
x"00",	-- Hex Addr	0C4A	3146
x"00",	-- Hex Addr	0C4B	3147
x"00",	-- Hex Addr	0C4C	3148
x"00",	-- Hex Addr	0C4D	3149
x"00",	-- Hex Addr	0C4E	3150
x"00",	-- Hex Addr	0C4F	3151
x"00",	-- Hex Addr	0C50	3152
x"00",	-- Hex Addr	0C51	3153
x"00",	-- Hex Addr	0C52	3154
x"00",	-- Hex Addr	0C53	3155
x"00",	-- Hex Addr	0C54	3156
x"00",	-- Hex Addr	0C55	3157
x"00",	-- Hex Addr	0C56	3158
x"00",	-- Hex Addr	0C57	3159
x"00",	-- Hex Addr	0C58	3160
x"00",	-- Hex Addr	0C59	3161
x"00",	-- Hex Addr	0C5A	3162
x"00",	-- Hex Addr	0C5B	3163
x"00",	-- Hex Addr	0C5C	3164
x"00",	-- Hex Addr	0C5D	3165
x"00",	-- Hex Addr	0C5E	3166
x"00",	-- Hex Addr	0C5F	3167
x"00",	-- Hex Addr	0C60	3168
x"00",	-- Hex Addr	0C61	3169
x"00",	-- Hex Addr	0C62	3170
x"00",	-- Hex Addr	0C63	3171
x"00",	-- Hex Addr	0C64	3172
x"00",	-- Hex Addr	0C65	3173
x"00",	-- Hex Addr	0C66	3174
x"00",	-- Hex Addr	0C67	3175
x"00",	-- Hex Addr	0C68	3176
x"00",	-- Hex Addr	0C69	3177
x"00",	-- Hex Addr	0C6A	3178
x"00",	-- Hex Addr	0C6B	3179
x"00",	-- Hex Addr	0C6C	3180
x"00",	-- Hex Addr	0C6D	3181
x"00",	-- Hex Addr	0C6E	3182
x"00",	-- Hex Addr	0C6F	3183
x"00",	-- Hex Addr	0C70	3184
x"00",	-- Hex Addr	0C71	3185
x"00",	-- Hex Addr	0C72	3186
x"00",	-- Hex Addr	0C73	3187
x"00",	-- Hex Addr	0C74	3188
x"00",	-- Hex Addr	0C75	3189
x"00",	-- Hex Addr	0C76	3190
x"00",	-- Hex Addr	0C77	3191
x"00",	-- Hex Addr	0C78	3192
x"00",	-- Hex Addr	0C79	3193
x"00",	-- Hex Addr	0C7A	3194
x"00",	-- Hex Addr	0C7B	3195
x"00",	-- Hex Addr	0C7C	3196
x"00",	-- Hex Addr	0C7D	3197
x"00",	-- Hex Addr	0C7E	3198
x"00",	-- Hex Addr	0C7F	3199
x"00",	-- Hex Addr	0C80	3200
x"00",	-- Hex Addr	0C81	3201
x"00",	-- Hex Addr	0C82	3202
x"00",	-- Hex Addr	0C83	3203
x"00",	-- Hex Addr	0C84	3204
x"00",	-- Hex Addr	0C85	3205
x"00",	-- Hex Addr	0C86	3206
x"00",	-- Hex Addr	0C87	3207
x"00",	-- Hex Addr	0C88	3208
x"00",	-- Hex Addr	0C89	3209
x"00",	-- Hex Addr	0C8A	3210
x"00",	-- Hex Addr	0C8B	3211
x"00",	-- Hex Addr	0C8C	3212
x"00",	-- Hex Addr	0C8D	3213
x"00",	-- Hex Addr	0C8E	3214
x"00",	-- Hex Addr	0C8F	3215
x"00",	-- Hex Addr	0C90	3216
x"00",	-- Hex Addr	0C91	3217
x"00",	-- Hex Addr	0C92	3218
x"00",	-- Hex Addr	0C93	3219
x"00",	-- Hex Addr	0C94	3220
x"00",	-- Hex Addr	0C95	3221
x"00",	-- Hex Addr	0C96	3222
x"00",	-- Hex Addr	0C97	3223
x"00",	-- Hex Addr	0C98	3224
x"00",	-- Hex Addr	0C99	3225
x"00",	-- Hex Addr	0C9A	3226
x"00",	-- Hex Addr	0C9B	3227
x"00",	-- Hex Addr	0C9C	3228
x"00",	-- Hex Addr	0C9D	3229
x"00",	-- Hex Addr	0C9E	3230
x"00",	-- Hex Addr	0C9F	3231
x"00",	-- Hex Addr	0CA0	3232
x"00",	-- Hex Addr	0CA1	3233
x"00",	-- Hex Addr	0CA2	3234
x"00",	-- Hex Addr	0CA3	3235
x"00",	-- Hex Addr	0CA4	3236
x"00",	-- Hex Addr	0CA5	3237
x"00",	-- Hex Addr	0CA6	3238
x"00",	-- Hex Addr	0CA7	3239
x"00",	-- Hex Addr	0CA8	3240
x"00",	-- Hex Addr	0CA9	3241
x"00",	-- Hex Addr	0CAA	3242
x"00",	-- Hex Addr	0CAB	3243
x"00",	-- Hex Addr	0CAC	3244
x"00",	-- Hex Addr	0CAD	3245
x"00",	-- Hex Addr	0CAE	3246
x"00",	-- Hex Addr	0CAF	3247
x"00",	-- Hex Addr	0CB0	3248
x"00",	-- Hex Addr	0CB1	3249
x"00",	-- Hex Addr	0CB2	3250
x"00",	-- Hex Addr	0CB3	3251
x"00",	-- Hex Addr	0CB4	3252
x"00",	-- Hex Addr	0CB5	3253
x"00",	-- Hex Addr	0CB6	3254
x"00",	-- Hex Addr	0CB7	3255
x"00",	-- Hex Addr	0CB8	3256
x"00",	-- Hex Addr	0CB9	3257
x"00",	-- Hex Addr	0CBA	3258
x"00",	-- Hex Addr	0CBB	3259
x"00",	-- Hex Addr	0CBC	3260
x"00",	-- Hex Addr	0CBD	3261
x"00",	-- Hex Addr	0CBE	3262
x"00",	-- Hex Addr	0CBF	3263
x"00",	-- Hex Addr	0CC0	3264
x"00",	-- Hex Addr	0CC1	3265
x"00",	-- Hex Addr	0CC2	3266
x"00",	-- Hex Addr	0CC3	3267
x"00",	-- Hex Addr	0CC4	3268
x"00",	-- Hex Addr	0CC5	3269
x"00",	-- Hex Addr	0CC6	3270
x"00",	-- Hex Addr	0CC7	3271
x"00",	-- Hex Addr	0CC8	3272
x"00",	-- Hex Addr	0CC9	3273
x"00",	-- Hex Addr	0CCA	3274
x"00",	-- Hex Addr	0CCB	3275
x"00",	-- Hex Addr	0CCC	3276
x"00",	-- Hex Addr	0CCD	3277
x"00",	-- Hex Addr	0CCE	3278
x"00",	-- Hex Addr	0CCF	3279
x"00",	-- Hex Addr	0CD0	3280
x"00",	-- Hex Addr	0CD1	3281
x"00",	-- Hex Addr	0CD2	3282
x"00",	-- Hex Addr	0CD3	3283
x"00",	-- Hex Addr	0CD4	3284
x"00",	-- Hex Addr	0CD5	3285
x"00",	-- Hex Addr	0CD6	3286
x"00",	-- Hex Addr	0CD7	3287
x"00",	-- Hex Addr	0CD8	3288
x"00",	-- Hex Addr	0CD9	3289
x"00",	-- Hex Addr	0CDA	3290
x"00",	-- Hex Addr	0CDB	3291
x"00",	-- Hex Addr	0CDC	3292
x"00",	-- Hex Addr	0CDD	3293
x"00",	-- Hex Addr	0CDE	3294
x"00",	-- Hex Addr	0CDF	3295
x"00",	-- Hex Addr	0CE0	3296
x"00",	-- Hex Addr	0CE1	3297
x"00",	-- Hex Addr	0CE2	3298
x"00",	-- Hex Addr	0CE3	3299
x"00",	-- Hex Addr	0CE4	3300
x"00",	-- Hex Addr	0CE5	3301
x"00",	-- Hex Addr	0CE6	3302
x"00",	-- Hex Addr	0CE7	3303
x"00",	-- Hex Addr	0CE8	3304
x"00",	-- Hex Addr	0CE9	3305
x"00",	-- Hex Addr	0CEA	3306
x"00",	-- Hex Addr	0CEB	3307
x"00",	-- Hex Addr	0CEC	3308
x"00",	-- Hex Addr	0CED	3309
x"00",	-- Hex Addr	0CEE	3310
x"00",	-- Hex Addr	0CEF	3311
x"00",	-- Hex Addr	0CF0	3312
x"00",	-- Hex Addr	0CF1	3313
x"00",	-- Hex Addr	0CF2	3314
x"00",	-- Hex Addr	0CF3	3315
x"00",	-- Hex Addr	0CF4	3316
x"00",	-- Hex Addr	0CF5	3317
x"00",	-- Hex Addr	0CF6	3318
x"00",	-- Hex Addr	0CF7	3319
x"00",	-- Hex Addr	0CF8	3320
x"00",	-- Hex Addr	0CF9	3321
x"00",	-- Hex Addr	0CFA	3322
x"00",	-- Hex Addr	0CFB	3323
x"00",	-- Hex Addr	0CFC	3324
x"00",	-- Hex Addr	0CFD	3325
x"00",	-- Hex Addr	0CFE	3326
x"00",	-- Hex Addr	0CFF	3327
x"00",	-- Hex Addr	0D00	3328
x"00",	-- Hex Addr	0D01	3329
x"00",	-- Hex Addr	0D02	3330
x"00",	-- Hex Addr	0D03	3331
x"00",	-- Hex Addr	0D04	3332
x"00",	-- Hex Addr	0D05	3333
x"00",	-- Hex Addr	0D06	3334
x"00",	-- Hex Addr	0D07	3335
x"00",	-- Hex Addr	0D08	3336
x"00",	-- Hex Addr	0D09	3337
x"00",	-- Hex Addr	0D0A	3338
x"00",	-- Hex Addr	0D0B	3339
x"00",	-- Hex Addr	0D0C	3340
x"00",	-- Hex Addr	0D0D	3341
x"00",	-- Hex Addr	0D0E	3342
x"00",	-- Hex Addr	0D0F	3343
x"00",	-- Hex Addr	0D10	3344
x"00",	-- Hex Addr	0D11	3345
x"00",	-- Hex Addr	0D12	3346
x"00",	-- Hex Addr	0D13	3347
x"00",	-- Hex Addr	0D14	3348
x"00",	-- Hex Addr	0D15	3349
x"00",	-- Hex Addr	0D16	3350
x"00",	-- Hex Addr	0D17	3351
x"00",	-- Hex Addr	0D18	3352
x"00",	-- Hex Addr	0D19	3353
x"00",	-- Hex Addr	0D1A	3354
x"00",	-- Hex Addr	0D1B	3355
x"00",	-- Hex Addr	0D1C	3356
x"00",	-- Hex Addr	0D1D	3357
x"00",	-- Hex Addr	0D1E	3358
x"00",	-- Hex Addr	0D1F	3359
x"00",	-- Hex Addr	0D20	3360
x"00",	-- Hex Addr	0D21	3361
x"00",	-- Hex Addr	0D22	3362
x"00",	-- Hex Addr	0D23	3363
x"00",	-- Hex Addr	0D24	3364
x"00",	-- Hex Addr	0D25	3365
x"00",	-- Hex Addr	0D26	3366
x"00",	-- Hex Addr	0D27	3367
x"00",	-- Hex Addr	0D28	3368
x"00",	-- Hex Addr	0D29	3369
x"00",	-- Hex Addr	0D2A	3370
x"00",	-- Hex Addr	0D2B	3371
x"00",	-- Hex Addr	0D2C	3372
x"00",	-- Hex Addr	0D2D	3373
x"00",	-- Hex Addr	0D2E	3374
x"00",	-- Hex Addr	0D2F	3375
x"00",	-- Hex Addr	0D30	3376
x"00",	-- Hex Addr	0D31	3377
x"00",	-- Hex Addr	0D32	3378
x"00",	-- Hex Addr	0D33	3379
x"00",	-- Hex Addr	0D34	3380
x"00",	-- Hex Addr	0D35	3381
x"00",	-- Hex Addr	0D36	3382
x"00",	-- Hex Addr	0D37	3383
x"00",	-- Hex Addr	0D38	3384
x"00",	-- Hex Addr	0D39	3385
x"00",	-- Hex Addr	0D3A	3386
x"00",	-- Hex Addr	0D3B	3387
x"00",	-- Hex Addr	0D3C	3388
x"00",	-- Hex Addr	0D3D	3389
x"00",	-- Hex Addr	0D3E	3390
x"00",	-- Hex Addr	0D3F	3391
x"00",	-- Hex Addr	0D40	3392
x"00",	-- Hex Addr	0D41	3393
x"00",	-- Hex Addr	0D42	3394
x"00",	-- Hex Addr	0D43	3395
x"00",	-- Hex Addr	0D44	3396
x"00",	-- Hex Addr	0D45	3397
x"00",	-- Hex Addr	0D46	3398
x"00",	-- Hex Addr	0D47	3399
x"00",	-- Hex Addr	0D48	3400
x"00",	-- Hex Addr	0D49	3401
x"00",	-- Hex Addr	0D4A	3402
x"00",	-- Hex Addr	0D4B	3403
x"00",	-- Hex Addr	0D4C	3404
x"00",	-- Hex Addr	0D4D	3405
x"00",	-- Hex Addr	0D4E	3406
x"00",	-- Hex Addr	0D4F	3407
x"00",	-- Hex Addr	0D50	3408
x"00",	-- Hex Addr	0D51	3409
x"00",	-- Hex Addr	0D52	3410
x"00",	-- Hex Addr	0D53	3411
x"00",	-- Hex Addr	0D54	3412
x"00",	-- Hex Addr	0D55	3413
x"00",	-- Hex Addr	0D56	3414
x"00",	-- Hex Addr	0D57	3415
x"00",	-- Hex Addr	0D58	3416
x"00",	-- Hex Addr	0D59	3417
x"00",	-- Hex Addr	0D5A	3418
x"00",	-- Hex Addr	0D5B	3419
x"00",	-- Hex Addr	0D5C	3420
x"00",	-- Hex Addr	0D5D	3421
x"00",	-- Hex Addr	0D5E	3422
x"00",	-- Hex Addr	0D5F	3423
x"00",	-- Hex Addr	0D60	3424
x"00",	-- Hex Addr	0D61	3425
x"00",	-- Hex Addr	0D62	3426
x"00",	-- Hex Addr	0D63	3427
x"00",	-- Hex Addr	0D64	3428
x"00",	-- Hex Addr	0D65	3429
x"00",	-- Hex Addr	0D66	3430
x"00",	-- Hex Addr	0D67	3431
x"00",	-- Hex Addr	0D68	3432
x"00",	-- Hex Addr	0D69	3433
x"00",	-- Hex Addr	0D6A	3434
x"00",	-- Hex Addr	0D6B	3435
x"00",	-- Hex Addr	0D6C	3436
x"00",	-- Hex Addr	0D6D	3437
x"00",	-- Hex Addr	0D6E	3438
x"00",	-- Hex Addr	0D6F	3439
x"00",	-- Hex Addr	0D70	3440
x"00",	-- Hex Addr	0D71	3441
x"00",	-- Hex Addr	0D72	3442
x"00",	-- Hex Addr	0D73	3443
x"00",	-- Hex Addr	0D74	3444
x"00",	-- Hex Addr	0D75	3445
x"00",	-- Hex Addr	0D76	3446
x"00",	-- Hex Addr	0D77	3447
x"00",	-- Hex Addr	0D78	3448
x"00",	-- Hex Addr	0D79	3449
x"00",	-- Hex Addr	0D7A	3450
x"00",	-- Hex Addr	0D7B	3451
x"00",	-- Hex Addr	0D7C	3452
x"00",	-- Hex Addr	0D7D	3453
x"00",	-- Hex Addr	0D7E	3454
x"00",	-- Hex Addr	0D7F	3455
x"00",	-- Hex Addr	0D80	3456
x"00",	-- Hex Addr	0D81	3457
x"00",	-- Hex Addr	0D82	3458
x"00",	-- Hex Addr	0D83	3459
x"00",	-- Hex Addr	0D84	3460
x"00",	-- Hex Addr	0D85	3461
x"00",	-- Hex Addr	0D86	3462
x"00",	-- Hex Addr	0D87	3463
x"00",	-- Hex Addr	0D88	3464
x"00",	-- Hex Addr	0D89	3465
x"00",	-- Hex Addr	0D8A	3466
x"00",	-- Hex Addr	0D8B	3467
x"00",	-- Hex Addr	0D8C	3468
x"00",	-- Hex Addr	0D8D	3469
x"00",	-- Hex Addr	0D8E	3470
x"00",	-- Hex Addr	0D8F	3471
x"00",	-- Hex Addr	0D90	3472
x"00",	-- Hex Addr	0D91	3473
x"00",	-- Hex Addr	0D92	3474
x"00",	-- Hex Addr	0D93	3475
x"00",	-- Hex Addr	0D94	3476
x"00",	-- Hex Addr	0D95	3477
x"00",	-- Hex Addr	0D96	3478
x"00",	-- Hex Addr	0D97	3479
x"00",	-- Hex Addr	0D98	3480
x"00",	-- Hex Addr	0D99	3481
x"00",	-- Hex Addr	0D9A	3482
x"00",	-- Hex Addr	0D9B	3483
x"00",	-- Hex Addr	0D9C	3484
x"00",	-- Hex Addr	0D9D	3485
x"00",	-- Hex Addr	0D9E	3486
x"00",	-- Hex Addr	0D9F	3487
x"00",	-- Hex Addr	0DA0	3488
x"00",	-- Hex Addr	0DA1	3489
x"00",	-- Hex Addr	0DA2	3490
x"00",	-- Hex Addr	0DA3	3491
x"00",	-- Hex Addr	0DA4	3492
x"00",	-- Hex Addr	0DA5	3493
x"00",	-- Hex Addr	0DA6	3494
x"00",	-- Hex Addr	0DA7	3495
x"00",	-- Hex Addr	0DA8	3496
x"00",	-- Hex Addr	0DA9	3497
x"00",	-- Hex Addr	0DAA	3498
x"00",	-- Hex Addr	0DAB	3499
x"00",	-- Hex Addr	0DAC	3500
x"00",	-- Hex Addr	0DAD	3501
x"00",	-- Hex Addr	0DAE	3502
x"00",	-- Hex Addr	0DAF	3503
x"00",	-- Hex Addr	0DB0	3504
x"00",	-- Hex Addr	0DB1	3505
x"00",	-- Hex Addr	0DB2	3506
x"00",	-- Hex Addr	0DB3	3507
x"00",	-- Hex Addr	0DB4	3508
x"00",	-- Hex Addr	0DB5	3509
x"00",	-- Hex Addr	0DB6	3510
x"00",	-- Hex Addr	0DB7	3511
x"00",	-- Hex Addr	0DB8	3512
x"00",	-- Hex Addr	0DB9	3513
x"00",	-- Hex Addr	0DBA	3514
x"00",	-- Hex Addr	0DBB	3515
x"00",	-- Hex Addr	0DBC	3516
x"00",	-- Hex Addr	0DBD	3517
x"00",	-- Hex Addr	0DBE	3518
x"00",	-- Hex Addr	0DBF	3519
x"00",	-- Hex Addr	0DC0	3520
x"00",	-- Hex Addr	0DC1	3521
x"00",	-- Hex Addr	0DC2	3522
x"00",	-- Hex Addr	0DC3	3523
x"00",	-- Hex Addr	0DC4	3524
x"00",	-- Hex Addr	0DC5	3525
x"00",	-- Hex Addr	0DC6	3526
x"00",	-- Hex Addr	0DC7	3527
x"00",	-- Hex Addr	0DC8	3528
x"00",	-- Hex Addr	0DC9	3529
x"00",	-- Hex Addr	0DCA	3530
x"00",	-- Hex Addr	0DCB	3531
x"00",	-- Hex Addr	0DCC	3532
x"00",	-- Hex Addr	0DCD	3533
x"00",	-- Hex Addr	0DCE	3534
x"00",	-- Hex Addr	0DCF	3535
x"00",	-- Hex Addr	0DD0	3536
x"00",	-- Hex Addr	0DD1	3537
x"00",	-- Hex Addr	0DD2	3538
x"00",	-- Hex Addr	0DD3	3539
x"00",	-- Hex Addr	0DD4	3540
x"00",	-- Hex Addr	0DD5	3541
x"00",	-- Hex Addr	0DD6	3542
x"00",	-- Hex Addr	0DD7	3543
x"00",	-- Hex Addr	0DD8	3544
x"00",	-- Hex Addr	0DD9	3545
x"00",	-- Hex Addr	0DDA	3546
x"00",	-- Hex Addr	0DDB	3547
x"00",	-- Hex Addr	0DDC	3548
x"00",	-- Hex Addr	0DDD	3549
x"00",	-- Hex Addr	0DDE	3550
x"00",	-- Hex Addr	0DDF	3551
x"00",	-- Hex Addr	0DE0	3552
x"00",	-- Hex Addr	0DE1	3553
x"00",	-- Hex Addr	0DE2	3554
x"00",	-- Hex Addr	0DE3	3555
x"00",	-- Hex Addr	0DE4	3556
x"00",	-- Hex Addr	0DE5	3557
x"00",	-- Hex Addr	0DE6	3558
x"00",	-- Hex Addr	0DE7	3559
x"00",	-- Hex Addr	0DE8	3560
x"00",	-- Hex Addr	0DE9	3561
x"00",	-- Hex Addr	0DEA	3562
x"00",	-- Hex Addr	0DEB	3563
x"00",	-- Hex Addr	0DEC	3564
x"00",	-- Hex Addr	0DED	3565
x"00",	-- Hex Addr	0DEE	3566
x"00",	-- Hex Addr	0DEF	3567
x"00",	-- Hex Addr	0DF0	3568
x"00",	-- Hex Addr	0DF1	3569
x"00",	-- Hex Addr	0DF2	3570
x"00",	-- Hex Addr	0DF3	3571
x"00",	-- Hex Addr	0DF4	3572
x"00",	-- Hex Addr	0DF5	3573
x"00",	-- Hex Addr	0DF6	3574
x"00",	-- Hex Addr	0DF7	3575
x"00",	-- Hex Addr	0DF8	3576
x"00",	-- Hex Addr	0DF9	3577
x"00",	-- Hex Addr	0DFA	3578
x"00",	-- Hex Addr	0DFB	3579
x"00",	-- Hex Addr	0DFC	3580
x"00",	-- Hex Addr	0DFD	3581
x"00",	-- Hex Addr	0DFE	3582
x"00",	-- Hex Addr	0DFF	3583
x"00",	-- Hex Addr	0E00	3584
x"00",	-- Hex Addr	0E01	3585
x"00",	-- Hex Addr	0E02	3586
x"00",	-- Hex Addr	0E03	3587
x"00",	-- Hex Addr	0E04	3588
x"00",	-- Hex Addr	0E05	3589
x"00",	-- Hex Addr	0E06	3590
x"00",	-- Hex Addr	0E07	3591
x"00",	-- Hex Addr	0E08	3592
x"00",	-- Hex Addr	0E09	3593
x"00",	-- Hex Addr	0E0A	3594
x"00",	-- Hex Addr	0E0B	3595
x"00",	-- Hex Addr	0E0C	3596
x"00",	-- Hex Addr	0E0D	3597
x"00",	-- Hex Addr	0E0E	3598
x"00",	-- Hex Addr	0E0F	3599
x"00",	-- Hex Addr	0E10	3600
x"00",	-- Hex Addr	0E11	3601
x"00",	-- Hex Addr	0E12	3602
x"00",	-- Hex Addr	0E13	3603
x"00",	-- Hex Addr	0E14	3604
x"00",	-- Hex Addr	0E15	3605
x"00",	-- Hex Addr	0E16	3606
x"00",	-- Hex Addr	0E17	3607
x"00",	-- Hex Addr	0E18	3608
x"00",	-- Hex Addr	0E19	3609
x"00",	-- Hex Addr	0E1A	3610
x"00",	-- Hex Addr	0E1B	3611
x"00",	-- Hex Addr	0E1C	3612
x"00",	-- Hex Addr	0E1D	3613
x"00",	-- Hex Addr	0E1E	3614
x"00",	-- Hex Addr	0E1F	3615
x"00",	-- Hex Addr	0E20	3616
x"00",	-- Hex Addr	0E21	3617
x"00",	-- Hex Addr	0E22	3618
x"00",	-- Hex Addr	0E23	3619
x"00",	-- Hex Addr	0E24	3620
x"00",	-- Hex Addr	0E25	3621
x"00",	-- Hex Addr	0E26	3622
x"00",	-- Hex Addr	0E27	3623
x"00",	-- Hex Addr	0E28	3624
x"00",	-- Hex Addr	0E29	3625
x"00",	-- Hex Addr	0E2A	3626
x"00",	-- Hex Addr	0E2B	3627
x"00",	-- Hex Addr	0E2C	3628
x"00",	-- Hex Addr	0E2D	3629
x"00",	-- Hex Addr	0E2E	3630
x"00",	-- Hex Addr	0E2F	3631
x"00",	-- Hex Addr	0E30	3632
x"00",	-- Hex Addr	0E31	3633
x"00",	-- Hex Addr	0E32	3634
x"00",	-- Hex Addr	0E33	3635
x"00",	-- Hex Addr	0E34	3636
x"00",	-- Hex Addr	0E35	3637
x"00",	-- Hex Addr	0E36	3638
x"00",	-- Hex Addr	0E37	3639
x"00",	-- Hex Addr	0E38	3640
x"00",	-- Hex Addr	0E39	3641
x"00",	-- Hex Addr	0E3A	3642
x"00",	-- Hex Addr	0E3B	3643
x"00",	-- Hex Addr	0E3C	3644
x"00",	-- Hex Addr	0E3D	3645
x"00",	-- Hex Addr	0E3E	3646
x"00",	-- Hex Addr	0E3F	3647
x"00",	-- Hex Addr	0E40	3648
x"00",	-- Hex Addr	0E41	3649
x"00",	-- Hex Addr	0E42	3650
x"00",	-- Hex Addr	0E43	3651
x"00",	-- Hex Addr	0E44	3652
x"00",	-- Hex Addr	0E45	3653
x"00",	-- Hex Addr	0E46	3654
x"00",	-- Hex Addr	0E47	3655
x"00",	-- Hex Addr	0E48	3656
x"00",	-- Hex Addr	0E49	3657
x"00",	-- Hex Addr	0E4A	3658
x"00",	-- Hex Addr	0E4B	3659
x"00",	-- Hex Addr	0E4C	3660
x"00",	-- Hex Addr	0E4D	3661
x"00",	-- Hex Addr	0E4E	3662
x"00",	-- Hex Addr	0E4F	3663
x"00",	-- Hex Addr	0E50	3664
x"00",	-- Hex Addr	0E51	3665
x"00",	-- Hex Addr	0E52	3666
x"00",	-- Hex Addr	0E53	3667
x"00",	-- Hex Addr	0E54	3668
x"00",	-- Hex Addr	0E55	3669
x"00",	-- Hex Addr	0E56	3670
x"00",	-- Hex Addr	0E57	3671
x"00",	-- Hex Addr	0E58	3672
x"00",	-- Hex Addr	0E59	3673
x"00",	-- Hex Addr	0E5A	3674
x"00",	-- Hex Addr	0E5B	3675
x"00",	-- Hex Addr	0E5C	3676
x"00",	-- Hex Addr	0E5D	3677
x"00",	-- Hex Addr	0E5E	3678
x"00",	-- Hex Addr	0E5F	3679
x"00",	-- Hex Addr	0E60	3680
x"00",	-- Hex Addr	0E61	3681
x"00",	-- Hex Addr	0E62	3682
x"00",	-- Hex Addr	0E63	3683
x"00",	-- Hex Addr	0E64	3684
x"00",	-- Hex Addr	0E65	3685
x"00",	-- Hex Addr	0E66	3686
x"00",	-- Hex Addr	0E67	3687
x"00",	-- Hex Addr	0E68	3688
x"00",	-- Hex Addr	0E69	3689
x"00",	-- Hex Addr	0E6A	3690
x"00",	-- Hex Addr	0E6B	3691
x"00",	-- Hex Addr	0E6C	3692
x"00",	-- Hex Addr	0E6D	3693
x"00",	-- Hex Addr	0E6E	3694
x"00",	-- Hex Addr	0E6F	3695
x"00",	-- Hex Addr	0E70	3696
x"00",	-- Hex Addr	0E71	3697
x"00",	-- Hex Addr	0E72	3698
x"00",	-- Hex Addr	0E73	3699
x"00",	-- Hex Addr	0E74	3700
x"00",	-- Hex Addr	0E75	3701
x"00",	-- Hex Addr	0E76	3702
x"00",	-- Hex Addr	0E77	3703
x"00",	-- Hex Addr	0E78	3704
x"00",	-- Hex Addr	0E79	3705
x"00",	-- Hex Addr	0E7A	3706
x"00",	-- Hex Addr	0E7B	3707
x"00",	-- Hex Addr	0E7C	3708
x"00",	-- Hex Addr	0E7D	3709
x"00",	-- Hex Addr	0E7E	3710
x"00",	-- Hex Addr	0E7F	3711
x"00",	-- Hex Addr	0E80	3712
x"00",	-- Hex Addr	0E81	3713
x"00",	-- Hex Addr	0E82	3714
x"00",	-- Hex Addr	0E83	3715
x"00",	-- Hex Addr	0E84	3716
x"00",	-- Hex Addr	0E85	3717
x"00",	-- Hex Addr	0E86	3718
x"00",	-- Hex Addr	0E87	3719
x"00",	-- Hex Addr	0E88	3720
x"00",	-- Hex Addr	0E89	3721
x"00",	-- Hex Addr	0E8A	3722
x"00",	-- Hex Addr	0E8B	3723
x"00",	-- Hex Addr	0E8C	3724
x"00",	-- Hex Addr	0E8D	3725
x"00",	-- Hex Addr	0E8E	3726
x"00",	-- Hex Addr	0E8F	3727
x"00",	-- Hex Addr	0E90	3728
x"00",	-- Hex Addr	0E91	3729
x"00",	-- Hex Addr	0E92	3730
x"00",	-- Hex Addr	0E93	3731
x"00",	-- Hex Addr	0E94	3732
x"00",	-- Hex Addr	0E95	3733
x"00",	-- Hex Addr	0E96	3734
x"00",	-- Hex Addr	0E97	3735
x"00",	-- Hex Addr	0E98	3736
x"00",	-- Hex Addr	0E99	3737
x"00",	-- Hex Addr	0E9A	3738
x"00",	-- Hex Addr	0E9B	3739
x"00",	-- Hex Addr	0E9C	3740
x"00",	-- Hex Addr	0E9D	3741
x"00",	-- Hex Addr	0E9E	3742
x"00",	-- Hex Addr	0E9F	3743
x"00",	-- Hex Addr	0EA0	3744
x"00",	-- Hex Addr	0EA1	3745
x"00",	-- Hex Addr	0EA2	3746
x"00",	-- Hex Addr	0EA3	3747
x"00",	-- Hex Addr	0EA4	3748
x"00",	-- Hex Addr	0EA5	3749
x"00",	-- Hex Addr	0EA6	3750
x"00",	-- Hex Addr	0EA7	3751
x"00",	-- Hex Addr	0EA8	3752
x"00",	-- Hex Addr	0EA9	3753
x"00",	-- Hex Addr	0EAA	3754
x"00",	-- Hex Addr	0EAB	3755
x"00",	-- Hex Addr	0EAC	3756
x"00",	-- Hex Addr	0EAD	3757
x"00",	-- Hex Addr	0EAE	3758
x"00",	-- Hex Addr	0EAF	3759
x"00",	-- Hex Addr	0EB0	3760
x"00",	-- Hex Addr	0EB1	3761
x"00",	-- Hex Addr	0EB2	3762
x"00",	-- Hex Addr	0EB3	3763
x"00",	-- Hex Addr	0EB4	3764
x"00",	-- Hex Addr	0EB5	3765
x"00",	-- Hex Addr	0EB6	3766
x"00",	-- Hex Addr	0EB7	3767
x"00",	-- Hex Addr	0EB8	3768
x"00",	-- Hex Addr	0EB9	3769
x"00",	-- Hex Addr	0EBA	3770
x"00",	-- Hex Addr	0EBB	3771
x"00",	-- Hex Addr	0EBC	3772
x"00",	-- Hex Addr	0EBD	3773
x"00",	-- Hex Addr	0EBE	3774
x"00",	-- Hex Addr	0EBF	3775
x"00",	-- Hex Addr	0EC0	3776
x"00",	-- Hex Addr	0EC1	3777
x"00",	-- Hex Addr	0EC2	3778
x"00",	-- Hex Addr	0EC3	3779
x"00",	-- Hex Addr	0EC4	3780
x"00",	-- Hex Addr	0EC5	3781
x"00",	-- Hex Addr	0EC6	3782
x"00",	-- Hex Addr	0EC7	3783
x"00",	-- Hex Addr	0EC8	3784
x"00",	-- Hex Addr	0EC9	3785
x"00",	-- Hex Addr	0ECA	3786
x"00",	-- Hex Addr	0ECB	3787
x"00",	-- Hex Addr	0ECC	3788
x"00",	-- Hex Addr	0ECD	3789
x"00",	-- Hex Addr	0ECE	3790
x"00",	-- Hex Addr	0ECF	3791
x"00",	-- Hex Addr	0ED0	3792
x"00",	-- Hex Addr	0ED1	3793
x"00",	-- Hex Addr	0ED2	3794
x"00",	-- Hex Addr	0ED3	3795
x"00",	-- Hex Addr	0ED4	3796
x"00",	-- Hex Addr	0ED5	3797
x"00",	-- Hex Addr	0ED6	3798
x"00",	-- Hex Addr	0ED7	3799
x"00",	-- Hex Addr	0ED8	3800
x"00",	-- Hex Addr	0ED9	3801
x"00",	-- Hex Addr	0EDA	3802
x"00",	-- Hex Addr	0EDB	3803
x"00",	-- Hex Addr	0EDC	3804
x"00",	-- Hex Addr	0EDD	3805
x"00",	-- Hex Addr	0EDE	3806
x"00",	-- Hex Addr	0EDF	3807
x"00",	-- Hex Addr	0EE0	3808
x"00",	-- Hex Addr	0EE1	3809
x"00",	-- Hex Addr	0EE2	3810
x"00",	-- Hex Addr	0EE3	3811
x"00",	-- Hex Addr	0EE4	3812
x"00",	-- Hex Addr	0EE5	3813
x"00",	-- Hex Addr	0EE6	3814
x"00",	-- Hex Addr	0EE7	3815
x"00",	-- Hex Addr	0EE8	3816
x"00",	-- Hex Addr	0EE9	3817
x"00",	-- Hex Addr	0EEA	3818
x"00",	-- Hex Addr	0EEB	3819
x"00",	-- Hex Addr	0EEC	3820
x"00",	-- Hex Addr	0EED	3821
x"00",	-- Hex Addr	0EEE	3822
x"00",	-- Hex Addr	0EEF	3823
x"00",	-- Hex Addr	0EF0	3824
x"00",	-- Hex Addr	0EF1	3825
x"00",	-- Hex Addr	0EF2	3826
x"00",	-- Hex Addr	0EF3	3827
x"00",	-- Hex Addr	0EF4	3828
x"00",	-- Hex Addr	0EF5	3829
x"00",	-- Hex Addr	0EF6	3830
x"00",	-- Hex Addr	0EF7	3831
x"00",	-- Hex Addr	0EF8	3832
x"00",	-- Hex Addr	0EF9	3833
x"00",	-- Hex Addr	0EFA	3834
x"00",	-- Hex Addr	0EFB	3835
x"00",	-- Hex Addr	0EFC	3836
x"00",	-- Hex Addr	0EFD	3837
x"00",	-- Hex Addr	0EFE	3838
x"00",	-- Hex Addr	0EFF	3839
x"00",	-- Hex Addr	0F00	3840
x"00",	-- Hex Addr	0F01	3841
x"00",	-- Hex Addr	0F02	3842
x"00",	-- Hex Addr	0F03	3843
x"00",	-- Hex Addr	0F04	3844
x"00",	-- Hex Addr	0F05	3845
x"00",	-- Hex Addr	0F06	3846
x"00",	-- Hex Addr	0F07	3847
x"00",	-- Hex Addr	0F08	3848
x"00",	-- Hex Addr	0F09	3849
x"00",	-- Hex Addr	0F0A	3850
x"00",	-- Hex Addr	0F0B	3851
x"00",	-- Hex Addr	0F0C	3852
x"00",	-- Hex Addr	0F0D	3853
x"00",	-- Hex Addr	0F0E	3854
x"00",	-- Hex Addr	0F0F	3855
x"00",	-- Hex Addr	0F10	3856
x"00",	-- Hex Addr	0F11	3857
x"00",	-- Hex Addr	0F12	3858
x"00",	-- Hex Addr	0F13	3859
x"00",	-- Hex Addr	0F14	3860
x"00",	-- Hex Addr	0F15	3861
x"00",	-- Hex Addr	0F16	3862
x"00",	-- Hex Addr	0F17	3863
x"00",	-- Hex Addr	0F18	3864
x"00",	-- Hex Addr	0F19	3865
x"00",	-- Hex Addr	0F1A	3866
x"00",	-- Hex Addr	0F1B	3867
x"00",	-- Hex Addr	0F1C	3868
x"00",	-- Hex Addr	0F1D	3869
x"00",	-- Hex Addr	0F1E	3870
x"00",	-- Hex Addr	0F1F	3871
x"00",	-- Hex Addr	0F20	3872
x"00",	-- Hex Addr	0F21	3873
x"00",	-- Hex Addr	0F22	3874
x"00",	-- Hex Addr	0F23	3875
x"00",	-- Hex Addr	0F24	3876
x"00",	-- Hex Addr	0F25	3877
x"00",	-- Hex Addr	0F26	3878
x"00",	-- Hex Addr	0F27	3879
x"00",	-- Hex Addr	0F28	3880
x"00",	-- Hex Addr	0F29	3881
x"00",	-- Hex Addr	0F2A	3882
x"00",	-- Hex Addr	0F2B	3883
x"00",	-- Hex Addr	0F2C	3884
x"00",	-- Hex Addr	0F2D	3885
x"00",	-- Hex Addr	0F2E	3886
x"00",	-- Hex Addr	0F2F	3887
x"00",	-- Hex Addr	0F30	3888
x"00",	-- Hex Addr	0F31	3889
x"00",	-- Hex Addr	0F32	3890
x"00",	-- Hex Addr	0F33	3891
x"00",	-- Hex Addr	0F34	3892
x"00",	-- Hex Addr	0F35	3893
x"00",	-- Hex Addr	0F36	3894
x"00",	-- Hex Addr	0F37	3895
x"00",	-- Hex Addr	0F38	3896
x"00",	-- Hex Addr	0F39	3897
x"00",	-- Hex Addr	0F3A	3898
x"00",	-- Hex Addr	0F3B	3899
x"00",	-- Hex Addr	0F3C	3900
x"00",	-- Hex Addr	0F3D	3901
x"00",	-- Hex Addr	0F3E	3902
x"00",	-- Hex Addr	0F3F	3903
x"00",	-- Hex Addr	0F40	3904
x"00",	-- Hex Addr	0F41	3905
x"00",	-- Hex Addr	0F42	3906
x"00",	-- Hex Addr	0F43	3907
x"00",	-- Hex Addr	0F44	3908
x"00",	-- Hex Addr	0F45	3909
x"00",	-- Hex Addr	0F46	3910
x"00",	-- Hex Addr	0F47	3911
x"00",	-- Hex Addr	0F48	3912
x"00",	-- Hex Addr	0F49	3913
x"00",	-- Hex Addr	0F4A	3914
x"00",	-- Hex Addr	0F4B	3915
x"00",	-- Hex Addr	0F4C	3916
x"00",	-- Hex Addr	0F4D	3917
x"00",	-- Hex Addr	0F4E	3918
x"00",	-- Hex Addr	0F4F	3919
x"00",	-- Hex Addr	0F50	3920
x"00",	-- Hex Addr	0F51	3921
x"00",	-- Hex Addr	0F52	3922
x"00",	-- Hex Addr	0F53	3923
x"00",	-- Hex Addr	0F54	3924
x"00",	-- Hex Addr	0F55	3925
x"00",	-- Hex Addr	0F56	3926
x"00",	-- Hex Addr	0F57	3927
x"00",	-- Hex Addr	0F58	3928
x"00",	-- Hex Addr	0F59	3929
x"00",	-- Hex Addr	0F5A	3930
x"00",	-- Hex Addr	0F5B	3931
x"00",	-- Hex Addr	0F5C	3932
x"00",	-- Hex Addr	0F5D	3933
x"00",	-- Hex Addr	0F5E	3934
x"00",	-- Hex Addr	0F5F	3935
x"00",	-- Hex Addr	0F60	3936
x"00",	-- Hex Addr	0F61	3937
x"00",	-- Hex Addr	0F62	3938
x"00",	-- Hex Addr	0F63	3939
x"00",	-- Hex Addr	0F64	3940
x"00",	-- Hex Addr	0F65	3941
x"00",	-- Hex Addr	0F66	3942
x"00",	-- Hex Addr	0F67	3943
x"00",	-- Hex Addr	0F68	3944
x"00",	-- Hex Addr	0F69	3945
x"00",	-- Hex Addr	0F6A	3946
x"00",	-- Hex Addr	0F6B	3947
x"00",	-- Hex Addr	0F6C	3948
x"00",	-- Hex Addr	0F6D	3949
x"00",	-- Hex Addr	0F6E	3950
x"00",	-- Hex Addr	0F6F	3951
x"00",	-- Hex Addr	0F70	3952
x"00",	-- Hex Addr	0F71	3953
x"00",	-- Hex Addr	0F72	3954
x"00",	-- Hex Addr	0F73	3955
x"00",	-- Hex Addr	0F74	3956
x"00",	-- Hex Addr	0F75	3957
x"00",	-- Hex Addr	0F76	3958
x"00",	-- Hex Addr	0F77	3959
x"00",	-- Hex Addr	0F78	3960
x"00",	-- Hex Addr	0F79	3961
x"00",	-- Hex Addr	0F7A	3962
x"00",	-- Hex Addr	0F7B	3963
x"00",	-- Hex Addr	0F7C	3964
x"00",	-- Hex Addr	0F7D	3965
x"00",	-- Hex Addr	0F7E	3966
x"00",	-- Hex Addr	0F7F	3967
x"00",	-- Hex Addr	0F80	3968
x"00",	-- Hex Addr	0F81	3969
x"00",	-- Hex Addr	0F82	3970
x"00",	-- Hex Addr	0F83	3971
x"00",	-- Hex Addr	0F84	3972
x"00",	-- Hex Addr	0F85	3973
x"00",	-- Hex Addr	0F86	3974
x"00",	-- Hex Addr	0F87	3975
x"00",	-- Hex Addr	0F88	3976
x"00",	-- Hex Addr	0F89	3977
x"00",	-- Hex Addr	0F8A	3978
x"00",	-- Hex Addr	0F8B	3979
x"00",	-- Hex Addr	0F8C	3980
x"00",	-- Hex Addr	0F8D	3981
x"00",	-- Hex Addr	0F8E	3982
x"00",	-- Hex Addr	0F8F	3983
x"00",	-- Hex Addr	0F90	3984
x"00",	-- Hex Addr	0F91	3985
x"00",	-- Hex Addr	0F92	3986
x"00",	-- Hex Addr	0F93	3987
x"00",	-- Hex Addr	0F94	3988
x"00",	-- Hex Addr	0F95	3989
x"00",	-- Hex Addr	0F96	3990
x"00",	-- Hex Addr	0F97	3991
x"00",	-- Hex Addr	0F98	3992
x"00",	-- Hex Addr	0F99	3993
x"00",	-- Hex Addr	0F9A	3994
x"00",	-- Hex Addr	0F9B	3995
x"00",	-- Hex Addr	0F9C	3996
x"00",	-- Hex Addr	0F9D	3997
x"00",	-- Hex Addr	0F9E	3998
x"00",	-- Hex Addr	0F9F	3999
x"00",	-- Hex Addr	0FA0	4000
x"00",	-- Hex Addr	0FA1	4001
x"00",	-- Hex Addr	0FA2	4002
x"00",	-- Hex Addr	0FA3	4003
x"00",	-- Hex Addr	0FA4	4004
x"00",	-- Hex Addr	0FA5	4005
x"00",	-- Hex Addr	0FA6	4006
x"00",	-- Hex Addr	0FA7	4007
x"00",	-- Hex Addr	0FA8	4008
x"00",	-- Hex Addr	0FA9	4009
x"00",	-- Hex Addr	0FAA	4010
x"00",	-- Hex Addr	0FAB	4011
x"00",	-- Hex Addr	0FAC	4012
x"00",	-- Hex Addr	0FAD	4013
x"00",	-- Hex Addr	0FAE	4014
x"00",	-- Hex Addr	0FAF	4015
x"00",	-- Hex Addr	0FB0	4016
x"00",	-- Hex Addr	0FB1	4017
x"00",	-- Hex Addr	0FB2	4018
x"00",	-- Hex Addr	0FB3	4019
x"00",	-- Hex Addr	0FB4	4020
x"00",	-- Hex Addr	0FB5	4021
x"00",	-- Hex Addr	0FB6	4022
x"00",	-- Hex Addr	0FB7	4023
x"00",	-- Hex Addr	0FB8	4024
x"00",	-- Hex Addr	0FB9	4025
x"00",	-- Hex Addr	0FBA	4026
x"00",	-- Hex Addr	0FBB	4027
x"00",	-- Hex Addr	0FBC	4028
x"00",	-- Hex Addr	0FBD	4029
x"00",	-- Hex Addr	0FBE	4030
x"00",	-- Hex Addr	0FBF	4031
x"00",	-- Hex Addr	0FC0	4032
x"00",	-- Hex Addr	0FC1	4033
x"00",	-- Hex Addr	0FC2	4034
x"00",	-- Hex Addr	0FC3	4035
x"00",	-- Hex Addr	0FC4	4036
x"00",	-- Hex Addr	0FC5	4037
x"00",	-- Hex Addr	0FC6	4038
x"00",	-- Hex Addr	0FC7	4039
x"00",	-- Hex Addr	0FC8	4040
x"00",	-- Hex Addr	0FC9	4041
x"00",	-- Hex Addr	0FCA	4042
x"00",	-- Hex Addr	0FCB	4043
x"00",	-- Hex Addr	0FCC	4044
x"00",	-- Hex Addr	0FCD	4045
x"00",	-- Hex Addr	0FCE	4046
x"00",	-- Hex Addr	0FCF	4047
x"00",	-- Hex Addr	0FD0	4048
x"00",	-- Hex Addr	0FD1	4049
x"00",	-- Hex Addr	0FD2	4050
x"00",	-- Hex Addr	0FD3	4051
x"00",	-- Hex Addr	0FD4	4052
x"00",	-- Hex Addr	0FD5	4053
x"00",	-- Hex Addr	0FD6	4054
x"00",	-- Hex Addr	0FD7	4055
x"00",	-- Hex Addr	0FD8	4056
x"00",	-- Hex Addr	0FD9	4057
x"00",	-- Hex Addr	0FDA	4058
x"00",	-- Hex Addr	0FDB	4059
x"00",	-- Hex Addr	0FDC	4060
x"00",	-- Hex Addr	0FDD	4061
x"00",	-- Hex Addr	0FDE	4062
x"00",	-- Hex Addr	0FDF	4063
x"00",	-- Hex Addr	0FE0	4064
x"00",	-- Hex Addr	0FE1	4065
x"00",	-- Hex Addr	0FE2	4066
x"00",	-- Hex Addr	0FE3	4067
x"00",	-- Hex Addr	0FE4	4068
x"00",	-- Hex Addr	0FE5	4069
x"00",	-- Hex Addr	0FE6	4070
x"00",	-- Hex Addr	0FE7	4071
x"00",	-- Hex Addr	0FE8	4072
x"00",	-- Hex Addr	0FE9	4073
x"00",	-- Hex Addr	0FEA	4074
x"00",	-- Hex Addr	0FEB	4075
x"00",	-- Hex Addr	0FEC	4076
x"00",	-- Hex Addr	0FED	4077
x"00",	-- Hex Addr	0FEE	4078
x"00",	-- Hex Addr	0FEF	4079
x"00",	-- Hex Addr	0FF0	4080
x"00",	-- Hex Addr	0FF1	4081
x"00",	-- Hex Addr	0FF2	4082
x"00",	-- Hex Addr	0FF3	4083
x"00",	-- Hex Addr	0FF4	4084
x"00",	-- Hex Addr	0FF5	4085
x"00",	-- Hex Addr	0FF6	4086
x"00",	-- Hex Addr	0FF7	4087
x"00",	-- Hex Addr	0FF8	4088
x"00",	-- Hex Addr	0FF9	4089
x"00",	-- Hex Addr	0FFA	4090
x"00",	-- Hex Addr	0FFB	4091
x"00",	-- Hex Addr	0FFC	4092
x"00",	-- Hex Addr	0FFD	4093
x"00",	-- Hex Addr	0FFE	4094
x"00",	-- Hex Addr	0FFF	4095
x"00",	-- Hex Addr	1000	4096
x"00",	-- Hex Addr	1001	4097
x"00",	-- Hex Addr	1002	4098
x"00",	-- Hex Addr	1003	4099
x"00",	-- Hex Addr	1004	4100
x"00",	-- Hex Addr	1005	4101
x"00",	-- Hex Addr	1006	4102
x"00",	-- Hex Addr	1007	4103
x"00",	-- Hex Addr	1008	4104
x"00",	-- Hex Addr	1009	4105
x"00",	-- Hex Addr	100A	4106
x"00",	-- Hex Addr	100B	4107
x"00",	-- Hex Addr	100C	4108
x"00",	-- Hex Addr	100D	4109
x"00",	-- Hex Addr	100E	4110
x"00",	-- Hex Addr	100F	4111
x"00",	-- Hex Addr	1010	4112
x"00",	-- Hex Addr	1011	4113
x"00",	-- Hex Addr	1012	4114
x"00",	-- Hex Addr	1013	4115
x"00",	-- Hex Addr	1014	4116
x"00",	-- Hex Addr	1015	4117
x"00",	-- Hex Addr	1016	4118
x"00",	-- Hex Addr	1017	4119
x"00",	-- Hex Addr	1018	4120
x"00",	-- Hex Addr	1019	4121
x"00",	-- Hex Addr	101A	4122
x"00",	-- Hex Addr	101B	4123
x"00",	-- Hex Addr	101C	4124
x"00",	-- Hex Addr	101D	4125
x"00",	-- Hex Addr	101E	4126
x"00",	-- Hex Addr	101F	4127
x"00",	-- Hex Addr	1020	4128
x"00",	-- Hex Addr	1021	4129
x"00",	-- Hex Addr	1022	4130
x"00",	-- Hex Addr	1023	4131
x"00",	-- Hex Addr	1024	4132
x"00",	-- Hex Addr	1025	4133
x"00",	-- Hex Addr	1026	4134
x"00",	-- Hex Addr	1027	4135
x"00",	-- Hex Addr	1028	4136
x"00",	-- Hex Addr	1029	4137
x"00",	-- Hex Addr	102A	4138
x"00",	-- Hex Addr	102B	4139
x"00",	-- Hex Addr	102C	4140
x"00",	-- Hex Addr	102D	4141
x"00",	-- Hex Addr	102E	4142
x"00",	-- Hex Addr	102F	4143
x"00",	-- Hex Addr	1030	4144
x"00",	-- Hex Addr	1031	4145
x"00",	-- Hex Addr	1032	4146
x"00",	-- Hex Addr	1033	4147
x"00",	-- Hex Addr	1034	4148
x"00",	-- Hex Addr	1035	4149
x"00",	-- Hex Addr	1036	4150
x"00",	-- Hex Addr	1037	4151
x"00",	-- Hex Addr	1038	4152
x"00",	-- Hex Addr	1039	4153
x"00",	-- Hex Addr	103A	4154
x"00",	-- Hex Addr	103B	4155
x"00",	-- Hex Addr	103C	4156
x"00",	-- Hex Addr	103D	4157
x"00",	-- Hex Addr	103E	4158
x"00",	-- Hex Addr	103F	4159
x"00",	-- Hex Addr	1040	4160
x"00",	-- Hex Addr	1041	4161
x"00",	-- Hex Addr	1042	4162
x"00",	-- Hex Addr	1043	4163
x"00",	-- Hex Addr	1044	4164
x"00",	-- Hex Addr	1045	4165
x"00",	-- Hex Addr	1046	4166
x"00",	-- Hex Addr	1047	4167
x"00",	-- Hex Addr	1048	4168
x"00",	-- Hex Addr	1049	4169
x"00",	-- Hex Addr	104A	4170
x"00",	-- Hex Addr	104B	4171
x"00",	-- Hex Addr	104C	4172
x"00",	-- Hex Addr	104D	4173
x"00",	-- Hex Addr	104E	4174
x"00",	-- Hex Addr	104F	4175
x"00",	-- Hex Addr	1050	4176
x"00",	-- Hex Addr	1051	4177
x"00",	-- Hex Addr	1052	4178
x"00",	-- Hex Addr	1053	4179
x"00",	-- Hex Addr	1054	4180
x"00",	-- Hex Addr	1055	4181
x"00",	-- Hex Addr	1056	4182
x"00",	-- Hex Addr	1057	4183
x"00",	-- Hex Addr	1058	4184
x"00",	-- Hex Addr	1059	4185
x"00",	-- Hex Addr	105A	4186
x"00",	-- Hex Addr	105B	4187
x"00",	-- Hex Addr	105C	4188
x"00",	-- Hex Addr	105D	4189
x"00",	-- Hex Addr	105E	4190
x"00",	-- Hex Addr	105F	4191
x"00",	-- Hex Addr	1060	4192
x"00",	-- Hex Addr	1061	4193
x"00",	-- Hex Addr	1062	4194
x"00",	-- Hex Addr	1063	4195
x"00",	-- Hex Addr	1064	4196
x"00",	-- Hex Addr	1065	4197
x"00",	-- Hex Addr	1066	4198
x"00",	-- Hex Addr	1067	4199
x"00",	-- Hex Addr	1068	4200
x"00",	-- Hex Addr	1069	4201
x"00",	-- Hex Addr	106A	4202
x"00",	-- Hex Addr	106B	4203
x"00",	-- Hex Addr	106C	4204
x"00",	-- Hex Addr	106D	4205
x"00",	-- Hex Addr	106E	4206
x"00",	-- Hex Addr	106F	4207
x"00",	-- Hex Addr	1070	4208
x"00",	-- Hex Addr	1071	4209
x"00",	-- Hex Addr	1072	4210
x"00",	-- Hex Addr	1073	4211
x"00",	-- Hex Addr	1074	4212
x"00",	-- Hex Addr	1075	4213
x"00",	-- Hex Addr	1076	4214
x"00",	-- Hex Addr	1077	4215
x"00",	-- Hex Addr	1078	4216
x"00",	-- Hex Addr	1079	4217
x"00",	-- Hex Addr	107A	4218
x"00",	-- Hex Addr	107B	4219
x"00",	-- Hex Addr	107C	4220
x"00",	-- Hex Addr	107D	4221
x"00",	-- Hex Addr	107E	4222
x"00",	-- Hex Addr	107F	4223
x"00",	-- Hex Addr	1080	4224
x"00",	-- Hex Addr	1081	4225
x"00",	-- Hex Addr	1082	4226
x"00",	-- Hex Addr	1083	4227
x"00",	-- Hex Addr	1084	4228
x"00",	-- Hex Addr	1085	4229
x"00",	-- Hex Addr	1086	4230
x"00",	-- Hex Addr	1087	4231
x"00",	-- Hex Addr	1088	4232
x"00",	-- Hex Addr	1089	4233
x"00",	-- Hex Addr	108A	4234
x"00",	-- Hex Addr	108B	4235
x"00",	-- Hex Addr	108C	4236
x"00",	-- Hex Addr	108D	4237
x"00",	-- Hex Addr	108E	4238
x"00",	-- Hex Addr	108F	4239
x"00",	-- Hex Addr	1090	4240
x"00",	-- Hex Addr	1091	4241
x"00",	-- Hex Addr	1092	4242
x"00",	-- Hex Addr	1093	4243
x"00",	-- Hex Addr	1094	4244
x"00",	-- Hex Addr	1095	4245
x"00",	-- Hex Addr	1096	4246
x"00",	-- Hex Addr	1097	4247
x"00",	-- Hex Addr	1098	4248
x"00",	-- Hex Addr	1099	4249
x"00",	-- Hex Addr	109A	4250
x"00",	-- Hex Addr	109B	4251
x"00",	-- Hex Addr	109C	4252
x"00",	-- Hex Addr	109D	4253
x"00",	-- Hex Addr	109E	4254
x"00",	-- Hex Addr	109F	4255
x"00",	-- Hex Addr	10A0	4256
x"00",	-- Hex Addr	10A1	4257
x"00",	-- Hex Addr	10A2	4258
x"00",	-- Hex Addr	10A3	4259
x"00",	-- Hex Addr	10A4	4260
x"00",	-- Hex Addr	10A5	4261
x"00",	-- Hex Addr	10A6	4262
x"00",	-- Hex Addr	10A7	4263
x"00",	-- Hex Addr	10A8	4264
x"00",	-- Hex Addr	10A9	4265
x"00",	-- Hex Addr	10AA	4266
x"00",	-- Hex Addr	10AB	4267
x"00",	-- Hex Addr	10AC	4268
x"00",	-- Hex Addr	10AD	4269
x"00",	-- Hex Addr	10AE	4270
x"00",	-- Hex Addr	10AF	4271
x"00",	-- Hex Addr	10B0	4272
x"00",	-- Hex Addr	10B1	4273
x"00",	-- Hex Addr	10B2	4274
x"00",	-- Hex Addr	10B3	4275
x"00",	-- Hex Addr	10B4	4276
x"00",	-- Hex Addr	10B5	4277
x"00",	-- Hex Addr	10B6	4278
x"00",	-- Hex Addr	10B7	4279
x"00",	-- Hex Addr	10B8	4280
x"00",	-- Hex Addr	10B9	4281
x"00",	-- Hex Addr	10BA	4282
x"00",	-- Hex Addr	10BB	4283
x"00",	-- Hex Addr	10BC	4284
x"00",	-- Hex Addr	10BD	4285
x"00",	-- Hex Addr	10BE	4286
x"00",	-- Hex Addr	10BF	4287
x"00",	-- Hex Addr	10C0	4288
x"00",	-- Hex Addr	10C1	4289
x"00",	-- Hex Addr	10C2	4290
x"00",	-- Hex Addr	10C3	4291
x"00",	-- Hex Addr	10C4	4292
x"00",	-- Hex Addr	10C5	4293
x"00",	-- Hex Addr	10C6	4294
x"00",	-- Hex Addr	10C7	4295
x"00",	-- Hex Addr	10C8	4296
x"00",	-- Hex Addr	10C9	4297
x"00",	-- Hex Addr	10CA	4298
x"00",	-- Hex Addr	10CB	4299
x"00",	-- Hex Addr	10CC	4300
x"00",	-- Hex Addr	10CD	4301
x"00",	-- Hex Addr	10CE	4302
x"00",	-- Hex Addr	10CF	4303
x"00",	-- Hex Addr	10D0	4304
x"00",	-- Hex Addr	10D1	4305
x"00",	-- Hex Addr	10D2	4306
x"00",	-- Hex Addr	10D3	4307
x"00",	-- Hex Addr	10D4	4308
x"00",	-- Hex Addr	10D5	4309
x"00",	-- Hex Addr	10D6	4310
x"00",	-- Hex Addr	10D7	4311
x"00",	-- Hex Addr	10D8	4312
x"00",	-- Hex Addr	10D9	4313
x"00",	-- Hex Addr	10DA	4314
x"00",	-- Hex Addr	10DB	4315
x"00",	-- Hex Addr	10DC	4316
x"00",	-- Hex Addr	10DD	4317
x"00",	-- Hex Addr	10DE	4318
x"00",	-- Hex Addr	10DF	4319
x"00",	-- Hex Addr	10E0	4320
x"00",	-- Hex Addr	10E1	4321
x"00",	-- Hex Addr	10E2	4322
x"00",	-- Hex Addr	10E3	4323
x"00",	-- Hex Addr	10E4	4324
x"00",	-- Hex Addr	10E5	4325
x"00",	-- Hex Addr	10E6	4326
x"00",	-- Hex Addr	10E7	4327
x"00",	-- Hex Addr	10E8	4328
x"00",	-- Hex Addr	10E9	4329
x"00",	-- Hex Addr	10EA	4330
x"00",	-- Hex Addr	10EB	4331
x"00",	-- Hex Addr	10EC	4332
x"00",	-- Hex Addr	10ED	4333
x"00",	-- Hex Addr	10EE	4334
x"00",	-- Hex Addr	10EF	4335
x"00",	-- Hex Addr	10F0	4336
x"00",	-- Hex Addr	10F1	4337
x"00",	-- Hex Addr	10F2	4338
x"00",	-- Hex Addr	10F3	4339
x"00",	-- Hex Addr	10F4	4340
x"00",	-- Hex Addr	10F5	4341
x"00",	-- Hex Addr	10F6	4342
x"00",	-- Hex Addr	10F7	4343
x"00",	-- Hex Addr	10F8	4344
x"00",	-- Hex Addr	10F9	4345
x"00",	-- Hex Addr	10FA	4346
x"00",	-- Hex Addr	10FB	4347
x"00",	-- Hex Addr	10FC	4348
x"00",	-- Hex Addr	10FD	4349
x"00",	-- Hex Addr	10FE	4350
x"00",	-- Hex Addr	10FF	4351
x"00",	-- Hex Addr	1100	4352
x"00",	-- Hex Addr	1101	4353
x"00",	-- Hex Addr	1102	4354
x"00",	-- Hex Addr	1103	4355
x"00",	-- Hex Addr	1104	4356
x"00",	-- Hex Addr	1105	4357
x"00",	-- Hex Addr	1106	4358
x"00",	-- Hex Addr	1107	4359
x"00",	-- Hex Addr	1108	4360
x"00",	-- Hex Addr	1109	4361
x"00",	-- Hex Addr	110A	4362
x"00",	-- Hex Addr	110B	4363
x"00",	-- Hex Addr	110C	4364
x"00",	-- Hex Addr	110D	4365
x"00",	-- Hex Addr	110E	4366
x"00",	-- Hex Addr	110F	4367
x"00",	-- Hex Addr	1110	4368
x"00",	-- Hex Addr	1111	4369
x"00",	-- Hex Addr	1112	4370
x"00",	-- Hex Addr	1113	4371
x"00",	-- Hex Addr	1114	4372
x"00",	-- Hex Addr	1115	4373
x"00",	-- Hex Addr	1116	4374
x"00",	-- Hex Addr	1117	4375
x"00",	-- Hex Addr	1118	4376
x"00",	-- Hex Addr	1119	4377
x"00",	-- Hex Addr	111A	4378
x"00",	-- Hex Addr	111B	4379
x"00",	-- Hex Addr	111C	4380
x"00",	-- Hex Addr	111D	4381
x"00",	-- Hex Addr	111E	4382
x"00",	-- Hex Addr	111F	4383
x"00",	-- Hex Addr	1120	4384
x"00",	-- Hex Addr	1121	4385
x"00",	-- Hex Addr	1122	4386
x"00",	-- Hex Addr	1123	4387
x"00",	-- Hex Addr	1124	4388
x"00",	-- Hex Addr	1125	4389
x"00",	-- Hex Addr	1126	4390
x"00",	-- Hex Addr	1127	4391
x"00",	-- Hex Addr	1128	4392
x"00",	-- Hex Addr	1129	4393
x"00",	-- Hex Addr	112A	4394
x"00",	-- Hex Addr	112B	4395
x"00",	-- Hex Addr	112C	4396
x"00",	-- Hex Addr	112D	4397
x"00",	-- Hex Addr	112E	4398
x"00",	-- Hex Addr	112F	4399
x"00",	-- Hex Addr	1130	4400
x"00",	-- Hex Addr	1131	4401
x"00",	-- Hex Addr	1132	4402
x"00",	-- Hex Addr	1133	4403
x"00",	-- Hex Addr	1134	4404
x"00",	-- Hex Addr	1135	4405
x"00",	-- Hex Addr	1136	4406
x"00",	-- Hex Addr	1137	4407
x"00",	-- Hex Addr	1138	4408
x"00",	-- Hex Addr	1139	4409
x"00",	-- Hex Addr	113A	4410
x"00",	-- Hex Addr	113B	4411
x"00",	-- Hex Addr	113C	4412
x"00",	-- Hex Addr	113D	4413
x"00",	-- Hex Addr	113E	4414
x"00",	-- Hex Addr	113F	4415
x"00",	-- Hex Addr	1140	4416
x"00",	-- Hex Addr	1141	4417
x"00",	-- Hex Addr	1142	4418
x"00",	-- Hex Addr	1143	4419
x"00",	-- Hex Addr	1144	4420
x"00",	-- Hex Addr	1145	4421
x"00",	-- Hex Addr	1146	4422
x"00",	-- Hex Addr	1147	4423
x"00",	-- Hex Addr	1148	4424
x"00",	-- Hex Addr	1149	4425
x"00",	-- Hex Addr	114A	4426
x"00",	-- Hex Addr	114B	4427
x"00",	-- Hex Addr	114C	4428
x"00",	-- Hex Addr	114D	4429
x"00",	-- Hex Addr	114E	4430
x"00",	-- Hex Addr	114F	4431
x"00",	-- Hex Addr	1150	4432
x"00",	-- Hex Addr	1151	4433
x"00",	-- Hex Addr	1152	4434
x"00",	-- Hex Addr	1153	4435
x"00",	-- Hex Addr	1154	4436
x"00",	-- Hex Addr	1155	4437
x"00",	-- Hex Addr	1156	4438
x"00",	-- Hex Addr	1157	4439
x"00",	-- Hex Addr	1158	4440
x"00",	-- Hex Addr	1159	4441
x"00",	-- Hex Addr	115A	4442
x"00",	-- Hex Addr	115B	4443
x"00",	-- Hex Addr	115C	4444
x"00",	-- Hex Addr	115D	4445
x"00",	-- Hex Addr	115E	4446
x"00",	-- Hex Addr	115F	4447
x"00",	-- Hex Addr	1160	4448
x"00",	-- Hex Addr	1161	4449
x"00",	-- Hex Addr	1162	4450
x"00",	-- Hex Addr	1163	4451
x"00",	-- Hex Addr	1164	4452
x"00",	-- Hex Addr	1165	4453
x"00",	-- Hex Addr	1166	4454
x"00",	-- Hex Addr	1167	4455
x"00",	-- Hex Addr	1168	4456
x"00",	-- Hex Addr	1169	4457
x"00",	-- Hex Addr	116A	4458
x"00",	-- Hex Addr	116B	4459
x"00",	-- Hex Addr	116C	4460
x"00",	-- Hex Addr	116D	4461
x"00",	-- Hex Addr	116E	4462
x"00",	-- Hex Addr	116F	4463
x"00",	-- Hex Addr	1170	4464
x"00",	-- Hex Addr	1171	4465
x"00",	-- Hex Addr	1172	4466
x"00",	-- Hex Addr	1173	4467
x"00",	-- Hex Addr	1174	4468
x"00",	-- Hex Addr	1175	4469
x"00",	-- Hex Addr	1176	4470
x"00",	-- Hex Addr	1177	4471
x"00",	-- Hex Addr	1178	4472
x"00",	-- Hex Addr	1179	4473
x"00",	-- Hex Addr	117A	4474
x"00",	-- Hex Addr	117B	4475
x"00",	-- Hex Addr	117C	4476
x"00",	-- Hex Addr	117D	4477
x"00",	-- Hex Addr	117E	4478
x"00",	-- Hex Addr	117F	4479
x"00",	-- Hex Addr	1180	4480
x"00",	-- Hex Addr	1181	4481
x"00",	-- Hex Addr	1182	4482
x"00",	-- Hex Addr	1183	4483
x"00",	-- Hex Addr	1184	4484
x"00",	-- Hex Addr	1185	4485
x"00",	-- Hex Addr	1186	4486
x"00",	-- Hex Addr	1187	4487
x"00",	-- Hex Addr	1188	4488
x"00",	-- Hex Addr	1189	4489
x"00",	-- Hex Addr	118A	4490
x"00",	-- Hex Addr	118B	4491
x"00",	-- Hex Addr	118C	4492
x"00",	-- Hex Addr	118D	4493
x"00",	-- Hex Addr	118E	4494
x"00",	-- Hex Addr	118F	4495
x"00",	-- Hex Addr	1190	4496
x"00",	-- Hex Addr	1191	4497
x"00",	-- Hex Addr	1192	4498
x"00",	-- Hex Addr	1193	4499
x"00",	-- Hex Addr	1194	4500
x"00",	-- Hex Addr	1195	4501
x"00",	-- Hex Addr	1196	4502
x"00",	-- Hex Addr	1197	4503
x"00",	-- Hex Addr	1198	4504
x"00",	-- Hex Addr	1199	4505
x"00",	-- Hex Addr	119A	4506
x"00",	-- Hex Addr	119B	4507
x"00",	-- Hex Addr	119C	4508
x"00",	-- Hex Addr	119D	4509
x"00",	-- Hex Addr	119E	4510
x"00",	-- Hex Addr	119F	4511
x"00",	-- Hex Addr	11A0	4512
x"00",	-- Hex Addr	11A1	4513
x"00",	-- Hex Addr	11A2	4514
x"00",	-- Hex Addr	11A3	4515
x"00",	-- Hex Addr	11A4	4516
x"00",	-- Hex Addr	11A5	4517
x"00",	-- Hex Addr	11A6	4518
x"00",	-- Hex Addr	11A7	4519
x"00",	-- Hex Addr	11A8	4520
x"00",	-- Hex Addr	11A9	4521
x"00",	-- Hex Addr	11AA	4522
x"00",	-- Hex Addr	11AB	4523
x"00",	-- Hex Addr	11AC	4524
x"00",	-- Hex Addr	11AD	4525
x"00",	-- Hex Addr	11AE	4526
x"00",	-- Hex Addr	11AF	4527
x"00",	-- Hex Addr	11B0	4528
x"00",	-- Hex Addr	11B1	4529
x"00",	-- Hex Addr	11B2	4530
x"00",	-- Hex Addr	11B3	4531
x"00",	-- Hex Addr	11B4	4532
x"00",	-- Hex Addr	11B5	4533
x"00",	-- Hex Addr	11B6	4534
x"00",	-- Hex Addr	11B7	4535
x"00",	-- Hex Addr	11B8	4536
x"00",	-- Hex Addr	11B9	4537
x"00",	-- Hex Addr	11BA	4538
x"00",	-- Hex Addr	11BB	4539
x"00",	-- Hex Addr	11BC	4540
x"00",	-- Hex Addr	11BD	4541
x"00",	-- Hex Addr	11BE	4542
x"00",	-- Hex Addr	11BF	4543
x"00",	-- Hex Addr	11C0	4544
x"00",	-- Hex Addr	11C1	4545
x"00",	-- Hex Addr	11C2	4546
x"00",	-- Hex Addr	11C3	4547
x"00",	-- Hex Addr	11C4	4548
x"00",	-- Hex Addr	11C5	4549
x"00",	-- Hex Addr	11C6	4550
x"00",	-- Hex Addr	11C7	4551
x"00",	-- Hex Addr	11C8	4552
x"00",	-- Hex Addr	11C9	4553
x"00",	-- Hex Addr	11CA	4554
x"00",	-- Hex Addr	11CB	4555
x"00",	-- Hex Addr	11CC	4556
x"00",	-- Hex Addr	11CD	4557
x"00",	-- Hex Addr	11CE	4558
x"00",	-- Hex Addr	11CF	4559
x"00",	-- Hex Addr	11D0	4560
x"00",	-- Hex Addr	11D1	4561
x"00",	-- Hex Addr	11D2	4562
x"00",	-- Hex Addr	11D3	4563
x"00",	-- Hex Addr	11D4	4564
x"00",	-- Hex Addr	11D5	4565
x"00",	-- Hex Addr	11D6	4566
x"00",	-- Hex Addr	11D7	4567
x"00",	-- Hex Addr	11D8	4568
x"00",	-- Hex Addr	11D9	4569
x"00",	-- Hex Addr	11DA	4570
x"00",	-- Hex Addr	11DB	4571
x"00",	-- Hex Addr	11DC	4572
x"00",	-- Hex Addr	11DD	4573
x"00",	-- Hex Addr	11DE	4574
x"00",	-- Hex Addr	11DF	4575
x"00",	-- Hex Addr	11E0	4576
x"00",	-- Hex Addr	11E1	4577
x"00",	-- Hex Addr	11E2	4578
x"00",	-- Hex Addr	11E3	4579
x"00",	-- Hex Addr	11E4	4580
x"00",	-- Hex Addr	11E5	4581
x"00",	-- Hex Addr	11E6	4582
x"00",	-- Hex Addr	11E7	4583
x"00",	-- Hex Addr	11E8	4584
x"00",	-- Hex Addr	11E9	4585
x"00",	-- Hex Addr	11EA	4586
x"00",	-- Hex Addr	11EB	4587
x"00",	-- Hex Addr	11EC	4588
x"00",	-- Hex Addr	11ED	4589
x"00",	-- Hex Addr	11EE	4590
x"00",	-- Hex Addr	11EF	4591
x"00",	-- Hex Addr	11F0	4592
x"00",	-- Hex Addr	11F1	4593
x"00",	-- Hex Addr	11F2	4594
x"00",	-- Hex Addr	11F3	4595
x"00",	-- Hex Addr	11F4	4596
x"00",	-- Hex Addr	11F5	4597
x"00",	-- Hex Addr	11F6	4598
x"00",	-- Hex Addr	11F7	4599
x"00",	-- Hex Addr	11F8	4600
x"00",	-- Hex Addr	11F9	4601
x"00",	-- Hex Addr	11FA	4602
x"00",	-- Hex Addr	11FB	4603
x"00",	-- Hex Addr	11FC	4604
x"00",	-- Hex Addr	11FD	4605
x"00",	-- Hex Addr	11FE	4606
x"00",	-- Hex Addr	11FF	4607
x"00",	-- Hex Addr	1200	4608
x"00",	-- Hex Addr	1201	4609
x"00",	-- Hex Addr	1202	4610
x"00",	-- Hex Addr	1203	4611
x"00",	-- Hex Addr	1204	4612
x"00",	-- Hex Addr	1205	4613
x"00",	-- Hex Addr	1206	4614
x"00",	-- Hex Addr	1207	4615
x"00",	-- Hex Addr	1208	4616
x"00",	-- Hex Addr	1209	4617
x"00",	-- Hex Addr	120A	4618
x"00",	-- Hex Addr	120B	4619
x"00",	-- Hex Addr	120C	4620
x"00",	-- Hex Addr	120D	4621
x"00",	-- Hex Addr	120E	4622
x"00",	-- Hex Addr	120F	4623
x"00",	-- Hex Addr	1210	4624
x"00",	-- Hex Addr	1211	4625
x"00",	-- Hex Addr	1212	4626
x"00",	-- Hex Addr	1213	4627
x"00",	-- Hex Addr	1214	4628
x"00",	-- Hex Addr	1215	4629
x"00",	-- Hex Addr	1216	4630
x"00",	-- Hex Addr	1217	4631
x"00",	-- Hex Addr	1218	4632
x"00",	-- Hex Addr	1219	4633
x"00",	-- Hex Addr	121A	4634
x"00",	-- Hex Addr	121B	4635
x"00",	-- Hex Addr	121C	4636
x"00",	-- Hex Addr	121D	4637
x"00",	-- Hex Addr	121E	4638
x"00",	-- Hex Addr	121F	4639
x"00",	-- Hex Addr	1220	4640
x"00",	-- Hex Addr	1221	4641
x"00",	-- Hex Addr	1222	4642
x"00",	-- Hex Addr	1223	4643
x"00",	-- Hex Addr	1224	4644
x"00",	-- Hex Addr	1225	4645
x"00",	-- Hex Addr	1226	4646
x"00",	-- Hex Addr	1227	4647
x"00",	-- Hex Addr	1228	4648
x"00",	-- Hex Addr	1229	4649
x"00",	-- Hex Addr	122A	4650
x"00",	-- Hex Addr	122B	4651
x"00",	-- Hex Addr	122C	4652
x"00",	-- Hex Addr	122D	4653
x"00",	-- Hex Addr	122E	4654
x"00",	-- Hex Addr	122F	4655
x"00",	-- Hex Addr	1230	4656
x"00",	-- Hex Addr	1231	4657
x"00",	-- Hex Addr	1232	4658
x"00",	-- Hex Addr	1233	4659
x"00",	-- Hex Addr	1234	4660
x"00",	-- Hex Addr	1235	4661
x"00",	-- Hex Addr	1236	4662
x"00",	-- Hex Addr	1237	4663
x"00",	-- Hex Addr	1238	4664
x"00",	-- Hex Addr	1239	4665
x"00",	-- Hex Addr	123A	4666
x"00",	-- Hex Addr	123B	4667
x"00",	-- Hex Addr	123C	4668
x"00",	-- Hex Addr	123D	4669
x"00",	-- Hex Addr	123E	4670
x"00",	-- Hex Addr	123F	4671
x"00",	-- Hex Addr	1240	4672
x"00",	-- Hex Addr	1241	4673
x"00",	-- Hex Addr	1242	4674
x"00",	-- Hex Addr	1243	4675
x"00",	-- Hex Addr	1244	4676
x"00",	-- Hex Addr	1245	4677
x"00",	-- Hex Addr	1246	4678
x"00",	-- Hex Addr	1247	4679
x"00",	-- Hex Addr	1248	4680
x"00",	-- Hex Addr	1249	4681
x"00",	-- Hex Addr	124A	4682
x"00",	-- Hex Addr	124B	4683
x"00",	-- Hex Addr	124C	4684
x"00",	-- Hex Addr	124D	4685
x"00",	-- Hex Addr	124E	4686
x"00",	-- Hex Addr	124F	4687
x"00",	-- Hex Addr	1250	4688
x"00",	-- Hex Addr	1251	4689
x"00",	-- Hex Addr	1252	4690
x"00",	-- Hex Addr	1253	4691
x"00",	-- Hex Addr	1254	4692
x"00",	-- Hex Addr	1255	4693
x"00",	-- Hex Addr	1256	4694
x"00",	-- Hex Addr	1257	4695
x"00",	-- Hex Addr	1258	4696
x"00",	-- Hex Addr	1259	4697
x"00",	-- Hex Addr	125A	4698
x"00",	-- Hex Addr	125B	4699
x"00",	-- Hex Addr	125C	4700
x"00",	-- Hex Addr	125D	4701
x"00",	-- Hex Addr	125E	4702
x"00",	-- Hex Addr	125F	4703
x"00",	-- Hex Addr	1260	4704
x"00",	-- Hex Addr	1261	4705
x"00",	-- Hex Addr	1262	4706
x"00",	-- Hex Addr	1263	4707
x"00",	-- Hex Addr	1264	4708
x"00",	-- Hex Addr	1265	4709
x"00",	-- Hex Addr	1266	4710
x"00",	-- Hex Addr	1267	4711
x"00",	-- Hex Addr	1268	4712
x"00",	-- Hex Addr	1269	4713
x"00",	-- Hex Addr	126A	4714
x"00",	-- Hex Addr	126B	4715
x"00",	-- Hex Addr	126C	4716
x"00",	-- Hex Addr	126D	4717
x"00",	-- Hex Addr	126E	4718
x"00",	-- Hex Addr	126F	4719
x"00",	-- Hex Addr	1270	4720
x"00",	-- Hex Addr	1271	4721
x"00",	-- Hex Addr	1272	4722
x"00",	-- Hex Addr	1273	4723
x"00",	-- Hex Addr	1274	4724
x"00",	-- Hex Addr	1275	4725
x"00",	-- Hex Addr	1276	4726
x"00",	-- Hex Addr	1277	4727
x"00",	-- Hex Addr	1278	4728
x"00",	-- Hex Addr	1279	4729
x"00",	-- Hex Addr	127A	4730
x"00",	-- Hex Addr	127B	4731
x"00",	-- Hex Addr	127C	4732
x"00",	-- Hex Addr	127D	4733
x"00",	-- Hex Addr	127E	4734
x"00",	-- Hex Addr	127F	4735
x"00",	-- Hex Addr	1280	4736
x"00",	-- Hex Addr	1281	4737
x"00",	-- Hex Addr	1282	4738
x"00",	-- Hex Addr	1283	4739
x"00",	-- Hex Addr	1284	4740
x"00",	-- Hex Addr	1285	4741
x"00",	-- Hex Addr	1286	4742
x"00",	-- Hex Addr	1287	4743
x"00",	-- Hex Addr	1288	4744
x"00",	-- Hex Addr	1289	4745
x"00",	-- Hex Addr	128A	4746
x"00",	-- Hex Addr	128B	4747
x"00",	-- Hex Addr	128C	4748
x"00",	-- Hex Addr	128D	4749
x"00",	-- Hex Addr	128E	4750
x"00",	-- Hex Addr	128F	4751
x"00",	-- Hex Addr	1290	4752
x"00",	-- Hex Addr	1291	4753
x"00",	-- Hex Addr	1292	4754
x"00",	-- Hex Addr	1293	4755
x"00",	-- Hex Addr	1294	4756
x"00",	-- Hex Addr	1295	4757
x"00",	-- Hex Addr	1296	4758
x"00",	-- Hex Addr	1297	4759
x"00",	-- Hex Addr	1298	4760
x"00",	-- Hex Addr	1299	4761
x"00",	-- Hex Addr	129A	4762
x"00",	-- Hex Addr	129B	4763
x"00",	-- Hex Addr	129C	4764
x"00",	-- Hex Addr	129D	4765
x"00",	-- Hex Addr	129E	4766
x"00",	-- Hex Addr	129F	4767
x"00",	-- Hex Addr	12A0	4768
x"00",	-- Hex Addr	12A1	4769
x"00",	-- Hex Addr	12A2	4770
x"00",	-- Hex Addr	12A3	4771
x"00",	-- Hex Addr	12A4	4772
x"00",	-- Hex Addr	12A5	4773
x"00",	-- Hex Addr	12A6	4774
x"00",	-- Hex Addr	12A7	4775
x"00",	-- Hex Addr	12A8	4776
x"00",	-- Hex Addr	12A9	4777
x"00",	-- Hex Addr	12AA	4778
x"00",	-- Hex Addr	12AB	4779
x"00",	-- Hex Addr	12AC	4780
x"00",	-- Hex Addr	12AD	4781
x"00",	-- Hex Addr	12AE	4782
x"00",	-- Hex Addr	12AF	4783
x"00",	-- Hex Addr	12B0	4784
x"00",	-- Hex Addr	12B1	4785
x"00",	-- Hex Addr	12B2	4786
x"00",	-- Hex Addr	12B3	4787
x"00",	-- Hex Addr	12B4	4788
x"00",	-- Hex Addr	12B5	4789
x"00",	-- Hex Addr	12B6	4790
x"00",	-- Hex Addr	12B7	4791
x"00",	-- Hex Addr	12B8	4792
x"00",	-- Hex Addr	12B9	4793
x"00",	-- Hex Addr	12BA	4794
x"00",	-- Hex Addr	12BB	4795
x"00",	-- Hex Addr	12BC	4796
x"00",	-- Hex Addr	12BD	4797
x"00",	-- Hex Addr	12BE	4798
x"00",	-- Hex Addr	12BF	4799
x"00",	-- Hex Addr	12C0	4800
x"00",	-- Hex Addr	12C1	4801
x"00",	-- Hex Addr	12C2	4802
x"00",	-- Hex Addr	12C3	4803
x"00",	-- Hex Addr	12C4	4804
x"00",	-- Hex Addr	12C5	4805
x"00",	-- Hex Addr	12C6	4806
x"00",	-- Hex Addr	12C7	4807
x"00",	-- Hex Addr	12C8	4808
x"00",	-- Hex Addr	12C9	4809
x"00",	-- Hex Addr	12CA	4810
x"00",	-- Hex Addr	12CB	4811
x"00",	-- Hex Addr	12CC	4812
x"00",	-- Hex Addr	12CD	4813
x"00",	-- Hex Addr	12CE	4814
x"00",	-- Hex Addr	12CF	4815
x"00",	-- Hex Addr	12D0	4816
x"00",	-- Hex Addr	12D1	4817
x"00",	-- Hex Addr	12D2	4818
x"00",	-- Hex Addr	12D3	4819
x"00",	-- Hex Addr	12D4	4820
x"00",	-- Hex Addr	12D5	4821
x"00",	-- Hex Addr	12D6	4822
x"00",	-- Hex Addr	12D7	4823
x"00",	-- Hex Addr	12D8	4824
x"00",	-- Hex Addr	12D9	4825
x"00",	-- Hex Addr	12DA	4826
x"00",	-- Hex Addr	12DB	4827
x"00",	-- Hex Addr	12DC	4828
x"00",	-- Hex Addr	12DD	4829
x"00",	-- Hex Addr	12DE	4830
x"00",	-- Hex Addr	12DF	4831
x"00",	-- Hex Addr	12E0	4832
x"00",	-- Hex Addr	12E1	4833
x"00",	-- Hex Addr	12E2	4834
x"00",	-- Hex Addr	12E3	4835
x"00",	-- Hex Addr	12E4	4836
x"00",	-- Hex Addr	12E5	4837
x"00",	-- Hex Addr	12E6	4838
x"00",	-- Hex Addr	12E7	4839
x"00",	-- Hex Addr	12E8	4840
x"00",	-- Hex Addr	12E9	4841
x"00",	-- Hex Addr	12EA	4842
x"00",	-- Hex Addr	12EB	4843
x"00",	-- Hex Addr	12EC	4844
x"00",	-- Hex Addr	12ED	4845
x"00",	-- Hex Addr	12EE	4846
x"00",	-- Hex Addr	12EF	4847
x"00",	-- Hex Addr	12F0	4848
x"00",	-- Hex Addr	12F1	4849
x"00",	-- Hex Addr	12F2	4850
x"00",	-- Hex Addr	12F3	4851
x"00",	-- Hex Addr	12F4	4852
x"00",	-- Hex Addr	12F5	4853
x"00",	-- Hex Addr	12F6	4854
x"00",	-- Hex Addr	12F7	4855
x"00",	-- Hex Addr	12F8	4856
x"00",	-- Hex Addr	12F9	4857
x"00",	-- Hex Addr	12FA	4858
x"00",	-- Hex Addr	12FB	4859
x"00",	-- Hex Addr	12FC	4860
x"00",	-- Hex Addr	12FD	4861
x"00",	-- Hex Addr	12FE	4862
x"00",	-- Hex Addr	12FF	4863
x"00",	-- Hex Addr	1300	4864
x"00",	-- Hex Addr	1301	4865
x"00",	-- Hex Addr	1302	4866
x"00",	-- Hex Addr	1303	4867
x"00",	-- Hex Addr	1304	4868
x"00",	-- Hex Addr	1305	4869
x"00",	-- Hex Addr	1306	4870
x"00",	-- Hex Addr	1307	4871
x"00",	-- Hex Addr	1308	4872
x"00",	-- Hex Addr	1309	4873
x"00",	-- Hex Addr	130A	4874
x"00",	-- Hex Addr	130B	4875
x"00",	-- Hex Addr	130C	4876
x"00",	-- Hex Addr	130D	4877
x"00",	-- Hex Addr	130E	4878
x"00",	-- Hex Addr	130F	4879
x"00",	-- Hex Addr	1310	4880
x"00",	-- Hex Addr	1311	4881
x"00",	-- Hex Addr	1312	4882
x"00",	-- Hex Addr	1313	4883
x"00",	-- Hex Addr	1314	4884
x"00",	-- Hex Addr	1315	4885
x"00",	-- Hex Addr	1316	4886
x"00",	-- Hex Addr	1317	4887
x"00",	-- Hex Addr	1318	4888
x"00",	-- Hex Addr	1319	4889
x"00",	-- Hex Addr	131A	4890
x"00",	-- Hex Addr	131B	4891
x"00",	-- Hex Addr	131C	4892
x"00",	-- Hex Addr	131D	4893
x"00",	-- Hex Addr	131E	4894
x"00",	-- Hex Addr	131F	4895
x"00",	-- Hex Addr	1320	4896
x"00",	-- Hex Addr	1321	4897
x"00",	-- Hex Addr	1322	4898
x"00",	-- Hex Addr	1323	4899
x"00",	-- Hex Addr	1324	4900
x"00",	-- Hex Addr	1325	4901
x"00",	-- Hex Addr	1326	4902
x"00",	-- Hex Addr	1327	4903
x"00",	-- Hex Addr	1328	4904
x"00",	-- Hex Addr	1329	4905
x"00",	-- Hex Addr	132A	4906
x"00",	-- Hex Addr	132B	4907
x"00",	-- Hex Addr	132C	4908
x"00",	-- Hex Addr	132D	4909
x"00",	-- Hex Addr	132E	4910
x"00",	-- Hex Addr	132F	4911
x"00",	-- Hex Addr	1330	4912
x"00",	-- Hex Addr	1331	4913
x"00",	-- Hex Addr	1332	4914
x"00",	-- Hex Addr	1333	4915
x"00",	-- Hex Addr	1334	4916
x"00",	-- Hex Addr	1335	4917
x"00",	-- Hex Addr	1336	4918
x"00",	-- Hex Addr	1337	4919
x"00",	-- Hex Addr	1338	4920
x"00",	-- Hex Addr	1339	4921
x"00",	-- Hex Addr	133A	4922
x"00",	-- Hex Addr	133B	4923
x"00",	-- Hex Addr	133C	4924
x"00",	-- Hex Addr	133D	4925
x"00",	-- Hex Addr	133E	4926
x"00",	-- Hex Addr	133F	4927
x"00",	-- Hex Addr	1340	4928
x"00",	-- Hex Addr	1341	4929
x"00",	-- Hex Addr	1342	4930
x"00",	-- Hex Addr	1343	4931
x"00",	-- Hex Addr	1344	4932
x"00",	-- Hex Addr	1345	4933
x"00",	-- Hex Addr	1346	4934
x"00",	-- Hex Addr	1347	4935
x"00",	-- Hex Addr	1348	4936
x"00",	-- Hex Addr	1349	4937
x"00",	-- Hex Addr	134A	4938
x"00",	-- Hex Addr	134B	4939
x"00",	-- Hex Addr	134C	4940
x"00",	-- Hex Addr	134D	4941
x"00",	-- Hex Addr	134E	4942
x"00",	-- Hex Addr	134F	4943
x"00",	-- Hex Addr	1350	4944
x"00",	-- Hex Addr	1351	4945
x"00",	-- Hex Addr	1352	4946
x"00",	-- Hex Addr	1353	4947
x"00",	-- Hex Addr	1354	4948
x"00",	-- Hex Addr	1355	4949
x"00",	-- Hex Addr	1356	4950
x"00",	-- Hex Addr	1357	4951
x"00",	-- Hex Addr	1358	4952
x"00",	-- Hex Addr	1359	4953
x"00",	-- Hex Addr	135A	4954
x"00",	-- Hex Addr	135B	4955
x"00",	-- Hex Addr	135C	4956
x"00",	-- Hex Addr	135D	4957
x"00",	-- Hex Addr	135E	4958
x"00",	-- Hex Addr	135F	4959
x"00",	-- Hex Addr	1360	4960
x"00",	-- Hex Addr	1361	4961
x"00",	-- Hex Addr	1362	4962
x"00",	-- Hex Addr	1363	4963
x"00",	-- Hex Addr	1364	4964
x"00",	-- Hex Addr	1365	4965
x"00",	-- Hex Addr	1366	4966
x"00",	-- Hex Addr	1367	4967
x"00",	-- Hex Addr	1368	4968
x"00",	-- Hex Addr	1369	4969
x"00",	-- Hex Addr	136A	4970
x"00",	-- Hex Addr	136B	4971
x"00",	-- Hex Addr	136C	4972
x"00",	-- Hex Addr	136D	4973
x"00",	-- Hex Addr	136E	4974
x"00",	-- Hex Addr	136F	4975
x"00",	-- Hex Addr	1370	4976
x"00",	-- Hex Addr	1371	4977
x"00",	-- Hex Addr	1372	4978
x"00",	-- Hex Addr	1373	4979
x"00",	-- Hex Addr	1374	4980
x"00",	-- Hex Addr	1375	4981
x"00",	-- Hex Addr	1376	4982
x"00",	-- Hex Addr	1377	4983
x"00",	-- Hex Addr	1378	4984
x"00",	-- Hex Addr	1379	4985
x"00",	-- Hex Addr	137A	4986
x"00",	-- Hex Addr	137B	4987
x"00",	-- Hex Addr	137C	4988
x"00",	-- Hex Addr	137D	4989
x"00",	-- Hex Addr	137E	4990
x"00",	-- Hex Addr	137F	4991
x"00",	-- Hex Addr	1380	4992
x"00",	-- Hex Addr	1381	4993
x"00",	-- Hex Addr	1382	4994
x"00",	-- Hex Addr	1383	4995
x"00",	-- Hex Addr	1384	4996
x"00",	-- Hex Addr	1385	4997
x"00",	-- Hex Addr	1386	4998
x"00",	-- Hex Addr	1387	4999
x"00",	-- Hex Addr	1388	5000
x"00",	-- Hex Addr	1389	5001
x"00",	-- Hex Addr	138A	5002
x"00",	-- Hex Addr	138B	5003
x"00",	-- Hex Addr	138C	5004
x"00",	-- Hex Addr	138D	5005
x"00",	-- Hex Addr	138E	5006
x"00",	-- Hex Addr	138F	5007
x"00",	-- Hex Addr	1390	5008
x"00",	-- Hex Addr	1391	5009
x"00",	-- Hex Addr	1392	5010
x"00",	-- Hex Addr	1393	5011
x"00",	-- Hex Addr	1394	5012
x"00",	-- Hex Addr	1395	5013
x"00",	-- Hex Addr	1396	5014
x"00",	-- Hex Addr	1397	5015
x"00",	-- Hex Addr	1398	5016
x"00",	-- Hex Addr	1399	5017
x"00",	-- Hex Addr	139A	5018
x"00",	-- Hex Addr	139B	5019
x"00",	-- Hex Addr	139C	5020
x"00",	-- Hex Addr	139D	5021
x"00",	-- Hex Addr	139E	5022
x"00",	-- Hex Addr	139F	5023
x"00",	-- Hex Addr	13A0	5024
x"00",	-- Hex Addr	13A1	5025
x"00",	-- Hex Addr	13A2	5026
x"00",	-- Hex Addr	13A3	5027
x"00",	-- Hex Addr	13A4	5028
x"00",	-- Hex Addr	13A5	5029
x"00",	-- Hex Addr	13A6	5030
x"00",	-- Hex Addr	13A7	5031
x"00",	-- Hex Addr	13A8	5032
x"00",	-- Hex Addr	13A9	5033
x"00",	-- Hex Addr	13AA	5034
x"00",	-- Hex Addr	13AB	5035
x"00",	-- Hex Addr	13AC	5036
x"00",	-- Hex Addr	13AD	5037
x"00",	-- Hex Addr	13AE	5038
x"00",	-- Hex Addr	13AF	5039
x"00",	-- Hex Addr	13B0	5040
x"00",	-- Hex Addr	13B1	5041
x"00",	-- Hex Addr	13B2	5042
x"00",	-- Hex Addr	13B3	5043
x"00",	-- Hex Addr	13B4	5044
x"00",	-- Hex Addr	13B5	5045
x"00",	-- Hex Addr	13B6	5046
x"00",	-- Hex Addr	13B7	5047
x"00",	-- Hex Addr	13B8	5048
x"00",	-- Hex Addr	13B9	5049
x"00",	-- Hex Addr	13BA	5050
x"00",	-- Hex Addr	13BB	5051
x"00",	-- Hex Addr	13BC	5052
x"00",	-- Hex Addr	13BD	5053
x"00",	-- Hex Addr	13BE	5054
x"00",	-- Hex Addr	13BF	5055
x"00",	-- Hex Addr	13C0	5056
x"00",	-- Hex Addr	13C1	5057
x"00",	-- Hex Addr	13C2	5058
x"00",	-- Hex Addr	13C3	5059
x"00",	-- Hex Addr	13C4	5060
x"00",	-- Hex Addr	13C5	5061
x"00",	-- Hex Addr	13C6	5062
x"00",	-- Hex Addr	13C7	5063
x"00",	-- Hex Addr	13C8	5064
x"00",	-- Hex Addr	13C9	5065
x"00",	-- Hex Addr	13CA	5066
x"00",	-- Hex Addr	13CB	5067
x"00",	-- Hex Addr	13CC	5068
x"00",	-- Hex Addr	13CD	5069
x"00",	-- Hex Addr	13CE	5070
x"00",	-- Hex Addr	13CF	5071
x"00",	-- Hex Addr	13D0	5072
x"00",	-- Hex Addr	13D1	5073
x"00",	-- Hex Addr	13D2	5074
x"00",	-- Hex Addr	13D3	5075
x"00",	-- Hex Addr	13D4	5076
x"00",	-- Hex Addr	13D5	5077
x"00",	-- Hex Addr	13D6	5078
x"00",	-- Hex Addr	13D7	5079
x"00",	-- Hex Addr	13D8	5080
x"00",	-- Hex Addr	13D9	5081
x"00",	-- Hex Addr	13DA	5082
x"00",	-- Hex Addr	13DB	5083
x"00",	-- Hex Addr	13DC	5084
x"00",	-- Hex Addr	13DD	5085
x"00",	-- Hex Addr	13DE	5086
x"00",	-- Hex Addr	13DF	5087
x"00",	-- Hex Addr	13E0	5088
x"00",	-- Hex Addr	13E1	5089
x"00",	-- Hex Addr	13E2	5090
x"00",	-- Hex Addr	13E3	5091
x"00",	-- Hex Addr	13E4	5092
x"00",	-- Hex Addr	13E5	5093
x"00",	-- Hex Addr	13E6	5094
x"00",	-- Hex Addr	13E7	5095
x"00",	-- Hex Addr	13E8	5096
x"00",	-- Hex Addr	13E9	5097
x"00",	-- Hex Addr	13EA	5098
x"00",	-- Hex Addr	13EB	5099
x"00",	-- Hex Addr	13EC	5100
x"00",	-- Hex Addr	13ED	5101
x"00",	-- Hex Addr	13EE	5102
x"00",	-- Hex Addr	13EF	5103
x"00",	-- Hex Addr	13F0	5104
x"00",	-- Hex Addr	13F1	5105
x"00",	-- Hex Addr	13F2	5106
x"00",	-- Hex Addr	13F3	5107
x"00",	-- Hex Addr	13F4	5108
x"00",	-- Hex Addr	13F5	5109
x"00",	-- Hex Addr	13F6	5110
x"00",	-- Hex Addr	13F7	5111
x"00",	-- Hex Addr	13F8	5112
x"00",	-- Hex Addr	13F9	5113
x"00",	-- Hex Addr	13FA	5114
x"00",	-- Hex Addr	13FB	5115
x"00",	-- Hex Addr	13FC	5116
x"00",	-- Hex Addr	13FD	5117
x"00",	-- Hex Addr	13FE	5118
x"00",	-- Hex Addr	13FF	5119
x"00",	-- Hex Addr	1400	5120
x"00",	-- Hex Addr	1401	5121
x"00",	-- Hex Addr	1402	5122
x"00",	-- Hex Addr	1403	5123
x"00",	-- Hex Addr	1404	5124
x"00",	-- Hex Addr	1405	5125
x"00",	-- Hex Addr	1406	5126
x"00",	-- Hex Addr	1407	5127
x"00",	-- Hex Addr	1408	5128
x"00",	-- Hex Addr	1409	5129
x"00",	-- Hex Addr	140A	5130
x"00",	-- Hex Addr	140B	5131
x"00",	-- Hex Addr	140C	5132
x"00",	-- Hex Addr	140D	5133
x"00",	-- Hex Addr	140E	5134
x"00",	-- Hex Addr	140F	5135
x"00",	-- Hex Addr	1410	5136
x"00",	-- Hex Addr	1411	5137
x"00",	-- Hex Addr	1412	5138
x"00",	-- Hex Addr	1413	5139
x"00",	-- Hex Addr	1414	5140
x"00",	-- Hex Addr	1415	5141
x"00",	-- Hex Addr	1416	5142
x"00",	-- Hex Addr	1417	5143
x"00",	-- Hex Addr	1418	5144
x"00",	-- Hex Addr	1419	5145
x"00",	-- Hex Addr	141A	5146
x"00",	-- Hex Addr	141B	5147
x"00",	-- Hex Addr	141C	5148
x"00",	-- Hex Addr	141D	5149
x"00",	-- Hex Addr	141E	5150
x"00",	-- Hex Addr	141F	5151
x"00",	-- Hex Addr	1420	5152
x"00",	-- Hex Addr	1421	5153
x"00",	-- Hex Addr	1422	5154
x"00",	-- Hex Addr	1423	5155
x"00",	-- Hex Addr	1424	5156
x"00",	-- Hex Addr	1425	5157
x"00",	-- Hex Addr	1426	5158
x"00",	-- Hex Addr	1427	5159
x"00",	-- Hex Addr	1428	5160
x"00",	-- Hex Addr	1429	5161
x"00",	-- Hex Addr	142A	5162
x"00",	-- Hex Addr	142B	5163
x"00",	-- Hex Addr	142C	5164
x"00",	-- Hex Addr	142D	5165
x"00",	-- Hex Addr	142E	5166
x"00",	-- Hex Addr	142F	5167
x"00",	-- Hex Addr	1430	5168
x"00",	-- Hex Addr	1431	5169
x"00",	-- Hex Addr	1432	5170
x"00",	-- Hex Addr	1433	5171
x"00",	-- Hex Addr	1434	5172
x"00",	-- Hex Addr	1435	5173
x"00",	-- Hex Addr	1436	5174
x"00",	-- Hex Addr	1437	5175
x"00",	-- Hex Addr	1438	5176
x"00",	-- Hex Addr	1439	5177
x"00",	-- Hex Addr	143A	5178
x"00",	-- Hex Addr	143B	5179
x"00",	-- Hex Addr	143C	5180
x"00",	-- Hex Addr	143D	5181
x"00",	-- Hex Addr	143E	5182
x"00",	-- Hex Addr	143F	5183
x"00",	-- Hex Addr	1440	5184
x"00",	-- Hex Addr	1441	5185
x"00",	-- Hex Addr	1442	5186
x"00",	-- Hex Addr	1443	5187
x"00",	-- Hex Addr	1444	5188
x"00",	-- Hex Addr	1445	5189
x"00",	-- Hex Addr	1446	5190
x"00",	-- Hex Addr	1447	5191
x"00",	-- Hex Addr	1448	5192
x"00",	-- Hex Addr	1449	5193
x"00",	-- Hex Addr	144A	5194
x"00",	-- Hex Addr	144B	5195
x"00",	-- Hex Addr	144C	5196
x"00",	-- Hex Addr	144D	5197
x"00",	-- Hex Addr	144E	5198
x"00",	-- Hex Addr	144F	5199
x"00",	-- Hex Addr	1450	5200
x"00",	-- Hex Addr	1451	5201
x"00",	-- Hex Addr	1452	5202
x"00",	-- Hex Addr	1453	5203
x"00",	-- Hex Addr	1454	5204
x"00",	-- Hex Addr	1455	5205
x"00",	-- Hex Addr	1456	5206
x"00",	-- Hex Addr	1457	5207
x"00",	-- Hex Addr	1458	5208
x"00",	-- Hex Addr	1459	5209
x"00",	-- Hex Addr	145A	5210
x"00",	-- Hex Addr	145B	5211
x"00",	-- Hex Addr	145C	5212
x"00",	-- Hex Addr	145D	5213
x"00",	-- Hex Addr	145E	5214
x"00",	-- Hex Addr	145F	5215
x"00",	-- Hex Addr	1460	5216
x"00",	-- Hex Addr	1461	5217
x"00",	-- Hex Addr	1462	5218
x"00",	-- Hex Addr	1463	5219
x"00",	-- Hex Addr	1464	5220
x"00",	-- Hex Addr	1465	5221
x"00",	-- Hex Addr	1466	5222
x"00",	-- Hex Addr	1467	5223
x"00",	-- Hex Addr	1468	5224
x"00",	-- Hex Addr	1469	5225
x"00",	-- Hex Addr	146A	5226
x"00",	-- Hex Addr	146B	5227
x"00",	-- Hex Addr	146C	5228
x"00",	-- Hex Addr	146D	5229
x"00",	-- Hex Addr	146E	5230
x"00",	-- Hex Addr	146F	5231
x"00",	-- Hex Addr	1470	5232
x"00",	-- Hex Addr	1471	5233
x"00",	-- Hex Addr	1472	5234
x"00",	-- Hex Addr	1473	5235
x"00",	-- Hex Addr	1474	5236
x"00",	-- Hex Addr	1475	5237
x"00",	-- Hex Addr	1476	5238
x"00",	-- Hex Addr	1477	5239
x"00",	-- Hex Addr	1478	5240
x"00",	-- Hex Addr	1479	5241
x"00",	-- Hex Addr	147A	5242
x"00",	-- Hex Addr	147B	5243
x"00",	-- Hex Addr	147C	5244
x"00",	-- Hex Addr	147D	5245
x"00",	-- Hex Addr	147E	5246
x"00",	-- Hex Addr	147F	5247
x"00",	-- Hex Addr	1480	5248
x"00",	-- Hex Addr	1481	5249
x"00",	-- Hex Addr	1482	5250
x"00",	-- Hex Addr	1483	5251
x"00",	-- Hex Addr	1484	5252
x"00",	-- Hex Addr	1485	5253
x"00",	-- Hex Addr	1486	5254
x"00",	-- Hex Addr	1487	5255
x"00",	-- Hex Addr	1488	5256
x"00",	-- Hex Addr	1489	5257
x"00",	-- Hex Addr	148A	5258
x"00",	-- Hex Addr	148B	5259
x"00",	-- Hex Addr	148C	5260
x"00",	-- Hex Addr	148D	5261
x"00",	-- Hex Addr	148E	5262
x"00",	-- Hex Addr	148F	5263
x"00",	-- Hex Addr	1490	5264
x"00",	-- Hex Addr	1491	5265
x"00",	-- Hex Addr	1492	5266
x"00",	-- Hex Addr	1493	5267
x"00",	-- Hex Addr	1494	5268
x"00",	-- Hex Addr	1495	5269
x"00",	-- Hex Addr	1496	5270
x"00",	-- Hex Addr	1497	5271
x"00",	-- Hex Addr	1498	5272
x"00",	-- Hex Addr	1499	5273
x"00",	-- Hex Addr	149A	5274
x"00",	-- Hex Addr	149B	5275
x"00",	-- Hex Addr	149C	5276
x"00",	-- Hex Addr	149D	5277
x"00",	-- Hex Addr	149E	5278
x"00",	-- Hex Addr	149F	5279
x"00",	-- Hex Addr	14A0	5280
x"00",	-- Hex Addr	14A1	5281
x"00",	-- Hex Addr	14A2	5282
x"00",	-- Hex Addr	14A3	5283
x"00",	-- Hex Addr	14A4	5284
x"00",	-- Hex Addr	14A5	5285
x"00",	-- Hex Addr	14A6	5286
x"00",	-- Hex Addr	14A7	5287
x"00",	-- Hex Addr	14A8	5288
x"00",	-- Hex Addr	14A9	5289
x"00",	-- Hex Addr	14AA	5290
x"00",	-- Hex Addr	14AB	5291
x"00",	-- Hex Addr	14AC	5292
x"00",	-- Hex Addr	14AD	5293
x"00",	-- Hex Addr	14AE	5294
x"00",	-- Hex Addr	14AF	5295
x"00",	-- Hex Addr	14B0	5296
x"00",	-- Hex Addr	14B1	5297
x"00",	-- Hex Addr	14B2	5298
x"00",	-- Hex Addr	14B3	5299
x"00",	-- Hex Addr	14B4	5300
x"00",	-- Hex Addr	14B5	5301
x"00",	-- Hex Addr	14B6	5302
x"00",	-- Hex Addr	14B7	5303
x"00",	-- Hex Addr	14B8	5304
x"00",	-- Hex Addr	14B9	5305
x"00",	-- Hex Addr	14BA	5306
x"00",	-- Hex Addr	14BB	5307
x"00",	-- Hex Addr	14BC	5308
x"00",	-- Hex Addr	14BD	5309
x"00",	-- Hex Addr	14BE	5310
x"00",	-- Hex Addr	14BF	5311
x"00",	-- Hex Addr	14C0	5312
x"00",	-- Hex Addr	14C1	5313
x"00",	-- Hex Addr	14C2	5314
x"00",	-- Hex Addr	14C3	5315
x"00",	-- Hex Addr	14C4	5316
x"00",	-- Hex Addr	14C5	5317
x"00",	-- Hex Addr	14C6	5318
x"00",	-- Hex Addr	14C7	5319
x"00",	-- Hex Addr	14C8	5320
x"00",	-- Hex Addr	14C9	5321
x"00",	-- Hex Addr	14CA	5322
x"00",	-- Hex Addr	14CB	5323
x"00",	-- Hex Addr	14CC	5324
x"00",	-- Hex Addr	14CD	5325
x"00",	-- Hex Addr	14CE	5326
x"00",	-- Hex Addr	14CF	5327
x"00",	-- Hex Addr	14D0	5328
x"00",	-- Hex Addr	14D1	5329
x"00",	-- Hex Addr	14D2	5330
x"00",	-- Hex Addr	14D3	5331
x"00",	-- Hex Addr	14D4	5332
x"00",	-- Hex Addr	14D5	5333
x"00",	-- Hex Addr	14D6	5334
x"00",	-- Hex Addr	14D7	5335
x"00",	-- Hex Addr	14D8	5336
x"00",	-- Hex Addr	14D9	5337
x"00",	-- Hex Addr	14DA	5338
x"00",	-- Hex Addr	14DB	5339
x"00",	-- Hex Addr	14DC	5340
x"00",	-- Hex Addr	14DD	5341
x"00",	-- Hex Addr	14DE	5342
x"00",	-- Hex Addr	14DF	5343
x"00",	-- Hex Addr	14E0	5344
x"00",	-- Hex Addr	14E1	5345
x"00",	-- Hex Addr	14E2	5346
x"00",	-- Hex Addr	14E3	5347
x"00",	-- Hex Addr	14E4	5348
x"00",	-- Hex Addr	14E5	5349
x"00",	-- Hex Addr	14E6	5350
x"00",	-- Hex Addr	14E7	5351
x"00",	-- Hex Addr	14E8	5352
x"00",	-- Hex Addr	14E9	5353
x"00",	-- Hex Addr	14EA	5354
x"00",	-- Hex Addr	14EB	5355
x"00",	-- Hex Addr	14EC	5356
x"00",	-- Hex Addr	14ED	5357
x"00",	-- Hex Addr	14EE	5358
x"00",	-- Hex Addr	14EF	5359
x"00",	-- Hex Addr	14F0	5360
x"00",	-- Hex Addr	14F1	5361
x"00",	-- Hex Addr	14F2	5362
x"00",	-- Hex Addr	14F3	5363
x"00",	-- Hex Addr	14F4	5364
x"00",	-- Hex Addr	14F5	5365
x"00",	-- Hex Addr	14F6	5366
x"00",	-- Hex Addr	14F7	5367
x"00",	-- Hex Addr	14F8	5368
x"00",	-- Hex Addr	14F9	5369
x"00",	-- Hex Addr	14FA	5370
x"00",	-- Hex Addr	14FB	5371
x"00",	-- Hex Addr	14FC	5372
x"00",	-- Hex Addr	14FD	5373
x"00",	-- Hex Addr	14FE	5374
x"00",	-- Hex Addr	14FF	5375
x"00",	-- Hex Addr	1500	5376
x"00",	-- Hex Addr	1501	5377
x"00",	-- Hex Addr	1502	5378
x"00",	-- Hex Addr	1503	5379
x"00",	-- Hex Addr	1504	5380
x"00",	-- Hex Addr	1505	5381
x"00",	-- Hex Addr	1506	5382
x"00",	-- Hex Addr	1507	5383
x"00",	-- Hex Addr	1508	5384
x"00",	-- Hex Addr	1509	5385
x"00",	-- Hex Addr	150A	5386
x"00",	-- Hex Addr	150B	5387
x"00",	-- Hex Addr	150C	5388
x"00",	-- Hex Addr	150D	5389
x"00",	-- Hex Addr	150E	5390
x"00",	-- Hex Addr	150F	5391
x"00",	-- Hex Addr	1510	5392
x"00",	-- Hex Addr	1511	5393
x"00",	-- Hex Addr	1512	5394
x"00",	-- Hex Addr	1513	5395
x"00",	-- Hex Addr	1514	5396
x"00",	-- Hex Addr	1515	5397
x"00",	-- Hex Addr	1516	5398
x"00",	-- Hex Addr	1517	5399
x"00",	-- Hex Addr	1518	5400
x"00",	-- Hex Addr	1519	5401
x"00",	-- Hex Addr	151A	5402
x"00",	-- Hex Addr	151B	5403
x"00",	-- Hex Addr	151C	5404
x"00",	-- Hex Addr	151D	5405
x"00",	-- Hex Addr	151E	5406
x"00",	-- Hex Addr	151F	5407
x"00",	-- Hex Addr	1520	5408
x"00",	-- Hex Addr	1521	5409
x"00",	-- Hex Addr	1522	5410
x"00",	-- Hex Addr	1523	5411
x"00",	-- Hex Addr	1524	5412
x"00",	-- Hex Addr	1525	5413
x"00",	-- Hex Addr	1526	5414
x"00",	-- Hex Addr	1527	5415
x"00",	-- Hex Addr	1528	5416
x"00",	-- Hex Addr	1529	5417
x"00",	-- Hex Addr	152A	5418
x"00",	-- Hex Addr	152B	5419
x"00",	-- Hex Addr	152C	5420
x"00",	-- Hex Addr	152D	5421
x"00",	-- Hex Addr	152E	5422
x"00",	-- Hex Addr	152F	5423
x"00",	-- Hex Addr	1530	5424
x"00",	-- Hex Addr	1531	5425
x"00",	-- Hex Addr	1532	5426
x"00",	-- Hex Addr	1533	5427
x"00",	-- Hex Addr	1534	5428
x"00",	-- Hex Addr	1535	5429
x"00",	-- Hex Addr	1536	5430
x"00",	-- Hex Addr	1537	5431
x"00",	-- Hex Addr	1538	5432
x"00",	-- Hex Addr	1539	5433
x"00",	-- Hex Addr	153A	5434
x"00",	-- Hex Addr	153B	5435
x"00",	-- Hex Addr	153C	5436
x"00",	-- Hex Addr	153D	5437
x"00",	-- Hex Addr	153E	5438
x"00",	-- Hex Addr	153F	5439
x"00",	-- Hex Addr	1540	5440
x"00",	-- Hex Addr	1541	5441
x"00",	-- Hex Addr	1542	5442
x"00",	-- Hex Addr	1543	5443
x"00",	-- Hex Addr	1544	5444
x"00",	-- Hex Addr	1545	5445
x"00",	-- Hex Addr	1546	5446
x"00",	-- Hex Addr	1547	5447
x"00",	-- Hex Addr	1548	5448
x"00",	-- Hex Addr	1549	5449
x"00",	-- Hex Addr	154A	5450
x"00",	-- Hex Addr	154B	5451
x"00",	-- Hex Addr	154C	5452
x"00",	-- Hex Addr	154D	5453
x"00",	-- Hex Addr	154E	5454
x"00",	-- Hex Addr	154F	5455
x"00",	-- Hex Addr	1550	5456
x"00",	-- Hex Addr	1551	5457
x"00",	-- Hex Addr	1552	5458
x"00",	-- Hex Addr	1553	5459
x"00",	-- Hex Addr	1554	5460
x"00",	-- Hex Addr	1555	5461
x"00",	-- Hex Addr	1556	5462
x"00",	-- Hex Addr	1557	5463
x"00",	-- Hex Addr	1558	5464
x"00",	-- Hex Addr	1559	5465
x"00",	-- Hex Addr	155A	5466
x"00",	-- Hex Addr	155B	5467
x"00",	-- Hex Addr	155C	5468
x"00",	-- Hex Addr	155D	5469
x"00",	-- Hex Addr	155E	5470
x"00",	-- Hex Addr	155F	5471
x"00",	-- Hex Addr	1560	5472
x"00",	-- Hex Addr	1561	5473
x"00",	-- Hex Addr	1562	5474
x"00",	-- Hex Addr	1563	5475
x"00",	-- Hex Addr	1564	5476
x"00",	-- Hex Addr	1565	5477
x"00",	-- Hex Addr	1566	5478
x"00",	-- Hex Addr	1567	5479
x"00",	-- Hex Addr	1568	5480
x"00",	-- Hex Addr	1569	5481
x"00",	-- Hex Addr	156A	5482
x"00",	-- Hex Addr	156B	5483
x"00",	-- Hex Addr	156C	5484
x"00",	-- Hex Addr	156D	5485
x"00",	-- Hex Addr	156E	5486
x"00",	-- Hex Addr	156F	5487
x"00",	-- Hex Addr	1570	5488
x"00",	-- Hex Addr	1571	5489
x"00",	-- Hex Addr	1572	5490
x"00",	-- Hex Addr	1573	5491
x"00",	-- Hex Addr	1574	5492
x"00",	-- Hex Addr	1575	5493
x"00",	-- Hex Addr	1576	5494
x"00",	-- Hex Addr	1577	5495
x"00",	-- Hex Addr	1578	5496
x"00",	-- Hex Addr	1579	5497
x"00",	-- Hex Addr	157A	5498
x"00",	-- Hex Addr	157B	5499
x"00",	-- Hex Addr	157C	5500
x"00",	-- Hex Addr	157D	5501
x"00",	-- Hex Addr	157E	5502
x"00",	-- Hex Addr	157F	5503
x"00",	-- Hex Addr	1580	5504
x"00",	-- Hex Addr	1581	5505
x"00",	-- Hex Addr	1582	5506
x"00",	-- Hex Addr	1583	5507
x"00",	-- Hex Addr	1584	5508
x"00",	-- Hex Addr	1585	5509
x"00",	-- Hex Addr	1586	5510
x"00",	-- Hex Addr	1587	5511
x"00",	-- Hex Addr	1588	5512
x"00",	-- Hex Addr	1589	5513
x"00",	-- Hex Addr	158A	5514
x"00",	-- Hex Addr	158B	5515
x"00",	-- Hex Addr	158C	5516
x"00",	-- Hex Addr	158D	5517
x"00",	-- Hex Addr	158E	5518
x"00",	-- Hex Addr	158F	5519
x"00",	-- Hex Addr	1590	5520
x"00",	-- Hex Addr	1591	5521
x"00",	-- Hex Addr	1592	5522
x"00",	-- Hex Addr	1593	5523
x"00",	-- Hex Addr	1594	5524
x"00",	-- Hex Addr	1595	5525
x"00",	-- Hex Addr	1596	5526
x"00",	-- Hex Addr	1597	5527
x"00",	-- Hex Addr	1598	5528
x"00",	-- Hex Addr	1599	5529
x"00",	-- Hex Addr	159A	5530
x"00",	-- Hex Addr	159B	5531
x"00",	-- Hex Addr	159C	5532
x"00",	-- Hex Addr	159D	5533
x"00",	-- Hex Addr	159E	5534
x"00",	-- Hex Addr	159F	5535
x"00",	-- Hex Addr	15A0	5536
x"00",	-- Hex Addr	15A1	5537
x"00",	-- Hex Addr	15A2	5538
x"00",	-- Hex Addr	15A3	5539
x"00",	-- Hex Addr	15A4	5540
x"00",	-- Hex Addr	15A5	5541
x"00",	-- Hex Addr	15A6	5542
x"00",	-- Hex Addr	15A7	5543
x"00",	-- Hex Addr	15A8	5544
x"00",	-- Hex Addr	15A9	5545
x"00",	-- Hex Addr	15AA	5546
x"00",	-- Hex Addr	15AB	5547
x"00",	-- Hex Addr	15AC	5548
x"00",	-- Hex Addr	15AD	5549
x"00",	-- Hex Addr	15AE	5550
x"00",	-- Hex Addr	15AF	5551
x"00",	-- Hex Addr	15B0	5552
x"00",	-- Hex Addr	15B1	5553
x"00",	-- Hex Addr	15B2	5554
x"00",	-- Hex Addr	15B3	5555
x"00",	-- Hex Addr	15B4	5556
x"00",	-- Hex Addr	15B5	5557
x"00",	-- Hex Addr	15B6	5558
x"00",	-- Hex Addr	15B7	5559
x"00",	-- Hex Addr	15B8	5560
x"00",	-- Hex Addr	15B9	5561
x"00",	-- Hex Addr	15BA	5562
x"00",	-- Hex Addr	15BB	5563
x"00",	-- Hex Addr	15BC	5564
x"00",	-- Hex Addr	15BD	5565
x"00",	-- Hex Addr	15BE	5566
x"00",	-- Hex Addr	15BF	5567
x"00",	-- Hex Addr	15C0	5568
x"00",	-- Hex Addr	15C1	5569
x"00",	-- Hex Addr	15C2	5570
x"00",	-- Hex Addr	15C3	5571
x"00",	-- Hex Addr	15C4	5572
x"00",	-- Hex Addr	15C5	5573
x"00",	-- Hex Addr	15C6	5574
x"00",	-- Hex Addr	15C7	5575
x"00",	-- Hex Addr	15C8	5576
x"00",	-- Hex Addr	15C9	5577
x"00",	-- Hex Addr	15CA	5578
x"00",	-- Hex Addr	15CB	5579
x"00",	-- Hex Addr	15CC	5580
x"00",	-- Hex Addr	15CD	5581
x"00",	-- Hex Addr	15CE	5582
x"00",	-- Hex Addr	15CF	5583
x"00",	-- Hex Addr	15D0	5584
x"00",	-- Hex Addr	15D1	5585
x"00",	-- Hex Addr	15D2	5586
x"00",	-- Hex Addr	15D3	5587
x"00",	-- Hex Addr	15D4	5588
x"00",	-- Hex Addr	15D5	5589
x"00",	-- Hex Addr	15D6	5590
x"00",	-- Hex Addr	15D7	5591
x"00",	-- Hex Addr	15D8	5592
x"00",	-- Hex Addr	15D9	5593
x"00",	-- Hex Addr	15DA	5594
x"00",	-- Hex Addr	15DB	5595
x"00",	-- Hex Addr	15DC	5596
x"00",	-- Hex Addr	15DD	5597
x"00",	-- Hex Addr	15DE	5598
x"00",	-- Hex Addr	15DF	5599
x"00",	-- Hex Addr	15E0	5600
x"00",	-- Hex Addr	15E1	5601
x"00",	-- Hex Addr	15E2	5602
x"00",	-- Hex Addr	15E3	5603
x"00",	-- Hex Addr	15E4	5604
x"00",	-- Hex Addr	15E5	5605
x"00",	-- Hex Addr	15E6	5606
x"00",	-- Hex Addr	15E7	5607
x"00",	-- Hex Addr	15E8	5608
x"00",	-- Hex Addr	15E9	5609
x"00",	-- Hex Addr	15EA	5610
x"00",	-- Hex Addr	15EB	5611
x"00",	-- Hex Addr	15EC	5612
x"00",	-- Hex Addr	15ED	5613
x"00",	-- Hex Addr	15EE	5614
x"00",	-- Hex Addr	15EF	5615
x"00",	-- Hex Addr	15F0	5616
x"00",	-- Hex Addr	15F1	5617
x"00",	-- Hex Addr	15F2	5618
x"00",	-- Hex Addr	15F3	5619
x"00",	-- Hex Addr	15F4	5620
x"00",	-- Hex Addr	15F5	5621
x"00",	-- Hex Addr	15F6	5622
x"00",	-- Hex Addr	15F7	5623
x"00",	-- Hex Addr	15F8	5624
x"00",	-- Hex Addr	15F9	5625
x"00",	-- Hex Addr	15FA	5626
x"00",	-- Hex Addr	15FB	5627
x"00",	-- Hex Addr	15FC	5628
x"00",	-- Hex Addr	15FD	5629
x"00",	-- Hex Addr	15FE	5630
x"00",	-- Hex Addr	15FF	5631
x"00",	-- Hex Addr	1600	5632
x"00",	-- Hex Addr	1601	5633
x"00",	-- Hex Addr	1602	5634
x"00",	-- Hex Addr	1603	5635
x"00",	-- Hex Addr	1604	5636
x"00",	-- Hex Addr	1605	5637
x"00",	-- Hex Addr	1606	5638
x"00",	-- Hex Addr	1607	5639
x"00",	-- Hex Addr	1608	5640
x"00",	-- Hex Addr	1609	5641
x"00",	-- Hex Addr	160A	5642
x"00",	-- Hex Addr	160B	5643
x"00",	-- Hex Addr	160C	5644
x"00",	-- Hex Addr	160D	5645
x"00",	-- Hex Addr	160E	5646
x"00",	-- Hex Addr	160F	5647
x"00",	-- Hex Addr	1610	5648
x"00",	-- Hex Addr	1611	5649
x"00",	-- Hex Addr	1612	5650
x"00",	-- Hex Addr	1613	5651
x"00",	-- Hex Addr	1614	5652
x"00",	-- Hex Addr	1615	5653
x"00",	-- Hex Addr	1616	5654
x"00",	-- Hex Addr	1617	5655
x"00",	-- Hex Addr	1618	5656
x"00",	-- Hex Addr	1619	5657
x"00",	-- Hex Addr	161A	5658
x"00",	-- Hex Addr	161B	5659
x"00",	-- Hex Addr	161C	5660
x"00",	-- Hex Addr	161D	5661
x"00",	-- Hex Addr	161E	5662
x"00",	-- Hex Addr	161F	5663
x"00",	-- Hex Addr	1620	5664
x"00",	-- Hex Addr	1621	5665
x"00",	-- Hex Addr	1622	5666
x"00",	-- Hex Addr	1623	5667
x"00",	-- Hex Addr	1624	5668
x"00",	-- Hex Addr	1625	5669
x"00",	-- Hex Addr	1626	5670
x"00",	-- Hex Addr	1627	5671
x"00",	-- Hex Addr	1628	5672
x"00",	-- Hex Addr	1629	5673
x"00",	-- Hex Addr	162A	5674
x"00",	-- Hex Addr	162B	5675
x"00",	-- Hex Addr	162C	5676
x"00",	-- Hex Addr	162D	5677
x"00",	-- Hex Addr	162E	5678
x"00",	-- Hex Addr	162F	5679
x"00",	-- Hex Addr	1630	5680
x"00",	-- Hex Addr	1631	5681
x"00",	-- Hex Addr	1632	5682
x"00",	-- Hex Addr	1633	5683
x"00",	-- Hex Addr	1634	5684
x"00",	-- Hex Addr	1635	5685
x"00",	-- Hex Addr	1636	5686
x"00",	-- Hex Addr	1637	5687
x"00",	-- Hex Addr	1638	5688
x"00",	-- Hex Addr	1639	5689
x"00",	-- Hex Addr	163A	5690
x"00",	-- Hex Addr	163B	5691
x"00",	-- Hex Addr	163C	5692
x"00",	-- Hex Addr	163D	5693
x"00",	-- Hex Addr	163E	5694
x"00",	-- Hex Addr	163F	5695
x"00",	-- Hex Addr	1640	5696
x"00",	-- Hex Addr	1641	5697
x"00",	-- Hex Addr	1642	5698
x"00",	-- Hex Addr	1643	5699
x"00",	-- Hex Addr	1644	5700
x"00",	-- Hex Addr	1645	5701
x"00",	-- Hex Addr	1646	5702
x"00",	-- Hex Addr	1647	5703
x"00",	-- Hex Addr	1648	5704
x"00",	-- Hex Addr	1649	5705
x"00",	-- Hex Addr	164A	5706
x"00",	-- Hex Addr	164B	5707
x"00",	-- Hex Addr	164C	5708
x"00",	-- Hex Addr	164D	5709
x"00",	-- Hex Addr	164E	5710
x"00",	-- Hex Addr	164F	5711
x"00",	-- Hex Addr	1650	5712
x"00",	-- Hex Addr	1651	5713
x"00",	-- Hex Addr	1652	5714
x"00",	-- Hex Addr	1653	5715
x"00",	-- Hex Addr	1654	5716
x"00",	-- Hex Addr	1655	5717
x"00",	-- Hex Addr	1656	5718
x"00",	-- Hex Addr	1657	5719
x"00",	-- Hex Addr	1658	5720
x"00",	-- Hex Addr	1659	5721
x"00",	-- Hex Addr	165A	5722
x"00",	-- Hex Addr	165B	5723
x"00",	-- Hex Addr	165C	5724
x"00",	-- Hex Addr	165D	5725
x"00",	-- Hex Addr	165E	5726
x"00",	-- Hex Addr	165F	5727
x"00",	-- Hex Addr	1660	5728
x"00",	-- Hex Addr	1661	5729
x"00",	-- Hex Addr	1662	5730
x"00",	-- Hex Addr	1663	5731
x"00",	-- Hex Addr	1664	5732
x"00",	-- Hex Addr	1665	5733
x"00",	-- Hex Addr	1666	5734
x"00",	-- Hex Addr	1667	5735
x"00",	-- Hex Addr	1668	5736
x"00",	-- Hex Addr	1669	5737
x"00",	-- Hex Addr	166A	5738
x"00",	-- Hex Addr	166B	5739
x"00",	-- Hex Addr	166C	5740
x"00",	-- Hex Addr	166D	5741
x"00",	-- Hex Addr	166E	5742
x"00",	-- Hex Addr	166F	5743
x"00",	-- Hex Addr	1670	5744
x"00",	-- Hex Addr	1671	5745
x"00",	-- Hex Addr	1672	5746
x"00",	-- Hex Addr	1673	5747
x"00",	-- Hex Addr	1674	5748
x"00",	-- Hex Addr	1675	5749
x"00",	-- Hex Addr	1676	5750
x"00",	-- Hex Addr	1677	5751
x"00",	-- Hex Addr	1678	5752
x"00",	-- Hex Addr	1679	5753
x"00",	-- Hex Addr	167A	5754
x"00",	-- Hex Addr	167B	5755
x"00",	-- Hex Addr	167C	5756
x"00",	-- Hex Addr	167D	5757
x"00",	-- Hex Addr	167E	5758
x"00",	-- Hex Addr	167F	5759
x"00",	-- Hex Addr	1680	5760
x"00",	-- Hex Addr	1681	5761
x"00",	-- Hex Addr	1682	5762
x"00",	-- Hex Addr	1683	5763
x"00",	-- Hex Addr	1684	5764
x"00",	-- Hex Addr	1685	5765
x"00",	-- Hex Addr	1686	5766
x"00",	-- Hex Addr	1687	5767
x"00",	-- Hex Addr	1688	5768
x"00",	-- Hex Addr	1689	5769
x"00",	-- Hex Addr	168A	5770
x"00",	-- Hex Addr	168B	5771
x"00",	-- Hex Addr	168C	5772
x"00",	-- Hex Addr	168D	5773
x"00",	-- Hex Addr	168E	5774
x"00",	-- Hex Addr	168F	5775
x"00",	-- Hex Addr	1690	5776
x"00",	-- Hex Addr	1691	5777
x"00",	-- Hex Addr	1692	5778
x"00",	-- Hex Addr	1693	5779
x"00",	-- Hex Addr	1694	5780
x"00",	-- Hex Addr	1695	5781
x"00",	-- Hex Addr	1696	5782
x"00",	-- Hex Addr	1697	5783
x"00",	-- Hex Addr	1698	5784
x"00",	-- Hex Addr	1699	5785
x"00",	-- Hex Addr	169A	5786
x"00",	-- Hex Addr	169B	5787
x"00",	-- Hex Addr	169C	5788
x"00",	-- Hex Addr	169D	5789
x"00",	-- Hex Addr	169E	5790
x"00",	-- Hex Addr	169F	5791
x"00",	-- Hex Addr	16A0	5792
x"00",	-- Hex Addr	16A1	5793
x"00",	-- Hex Addr	16A2	5794
x"00",	-- Hex Addr	16A3	5795
x"00",	-- Hex Addr	16A4	5796
x"00",	-- Hex Addr	16A5	5797
x"00",	-- Hex Addr	16A6	5798
x"00",	-- Hex Addr	16A7	5799
x"00",	-- Hex Addr	16A8	5800
x"00",	-- Hex Addr	16A9	5801
x"00",	-- Hex Addr	16AA	5802
x"00",	-- Hex Addr	16AB	5803
x"00",	-- Hex Addr	16AC	5804
x"00",	-- Hex Addr	16AD	5805
x"00",	-- Hex Addr	16AE	5806
x"00",	-- Hex Addr	16AF	5807
x"00",	-- Hex Addr	16B0	5808
x"00",	-- Hex Addr	16B1	5809
x"00",	-- Hex Addr	16B2	5810
x"00",	-- Hex Addr	16B3	5811
x"00",	-- Hex Addr	16B4	5812
x"00",	-- Hex Addr	16B5	5813
x"00",	-- Hex Addr	16B6	5814
x"00",	-- Hex Addr	16B7	5815
x"00",	-- Hex Addr	16B8	5816
x"00",	-- Hex Addr	16B9	5817
x"00",	-- Hex Addr	16BA	5818
x"00",	-- Hex Addr	16BB	5819
x"00",	-- Hex Addr	16BC	5820
x"00",	-- Hex Addr	16BD	5821
x"00",	-- Hex Addr	16BE	5822
x"00",	-- Hex Addr	16BF	5823
x"00",	-- Hex Addr	16C0	5824
x"00",	-- Hex Addr	16C1	5825
x"00",	-- Hex Addr	16C2	5826
x"00",	-- Hex Addr	16C3	5827
x"00",	-- Hex Addr	16C4	5828
x"00",	-- Hex Addr	16C5	5829
x"00",	-- Hex Addr	16C6	5830
x"00",	-- Hex Addr	16C7	5831
x"00",	-- Hex Addr	16C8	5832
x"00",	-- Hex Addr	16C9	5833
x"00",	-- Hex Addr	16CA	5834
x"00",	-- Hex Addr	16CB	5835
x"00",	-- Hex Addr	16CC	5836
x"00",	-- Hex Addr	16CD	5837
x"00",	-- Hex Addr	16CE	5838
x"00",	-- Hex Addr	16CF	5839
x"00",	-- Hex Addr	16D0	5840
x"00",	-- Hex Addr	16D1	5841
x"00",	-- Hex Addr	16D2	5842
x"00",	-- Hex Addr	16D3	5843
x"00",	-- Hex Addr	16D4	5844
x"00",	-- Hex Addr	16D5	5845
x"00",	-- Hex Addr	16D6	5846
x"00",	-- Hex Addr	16D7	5847
x"00",	-- Hex Addr	16D8	5848
x"00",	-- Hex Addr	16D9	5849
x"00",	-- Hex Addr	16DA	5850
x"00",	-- Hex Addr	16DB	5851
x"00",	-- Hex Addr	16DC	5852
x"00",	-- Hex Addr	16DD	5853
x"00",	-- Hex Addr	16DE	5854
x"00",	-- Hex Addr	16DF	5855
x"00",	-- Hex Addr	16E0	5856
x"00",	-- Hex Addr	16E1	5857
x"00",	-- Hex Addr	16E2	5858
x"00",	-- Hex Addr	16E3	5859
x"00",	-- Hex Addr	16E4	5860
x"00",	-- Hex Addr	16E5	5861
x"00",	-- Hex Addr	16E6	5862
x"00",	-- Hex Addr	16E7	5863
x"00",	-- Hex Addr	16E8	5864
x"00",	-- Hex Addr	16E9	5865
x"00",	-- Hex Addr	16EA	5866
x"00",	-- Hex Addr	16EB	5867
x"00",	-- Hex Addr	16EC	5868
x"00",	-- Hex Addr	16ED	5869
x"00",	-- Hex Addr	16EE	5870
x"00",	-- Hex Addr	16EF	5871
x"00",	-- Hex Addr	16F0	5872
x"00",	-- Hex Addr	16F1	5873
x"00",	-- Hex Addr	16F2	5874
x"00",	-- Hex Addr	16F3	5875
x"00",	-- Hex Addr	16F4	5876
x"00",	-- Hex Addr	16F5	5877
x"00",	-- Hex Addr	16F6	5878
x"00",	-- Hex Addr	16F7	5879
x"00",	-- Hex Addr	16F8	5880
x"00",	-- Hex Addr	16F9	5881
x"00",	-- Hex Addr	16FA	5882
x"00",	-- Hex Addr	16FB	5883
x"00",	-- Hex Addr	16FC	5884
x"00",	-- Hex Addr	16FD	5885
x"00",	-- Hex Addr	16FE	5886
x"00",	-- Hex Addr	16FF	5887
x"00",	-- Hex Addr	1700	5888
x"00",	-- Hex Addr	1701	5889
x"00",	-- Hex Addr	1702	5890
x"00",	-- Hex Addr	1703	5891
x"00",	-- Hex Addr	1704	5892
x"00",	-- Hex Addr	1705	5893
x"00",	-- Hex Addr	1706	5894
x"00",	-- Hex Addr	1707	5895
x"00",	-- Hex Addr	1708	5896
x"00",	-- Hex Addr	1709	5897
x"00",	-- Hex Addr	170A	5898
x"00",	-- Hex Addr	170B	5899
x"00",	-- Hex Addr	170C	5900
x"00",	-- Hex Addr	170D	5901
x"00",	-- Hex Addr	170E	5902
x"00",	-- Hex Addr	170F	5903
x"00",	-- Hex Addr	1710	5904
x"00",	-- Hex Addr	1711	5905
x"00",	-- Hex Addr	1712	5906
x"00",	-- Hex Addr	1713	5907
x"00",	-- Hex Addr	1714	5908
x"00",	-- Hex Addr	1715	5909
x"00",	-- Hex Addr	1716	5910
x"00",	-- Hex Addr	1717	5911
x"00",	-- Hex Addr	1718	5912
x"00",	-- Hex Addr	1719	5913
x"00",	-- Hex Addr	171A	5914
x"00",	-- Hex Addr	171B	5915
x"00",	-- Hex Addr	171C	5916
x"00",	-- Hex Addr	171D	5917
x"00",	-- Hex Addr	171E	5918
x"00",	-- Hex Addr	171F	5919
x"00",	-- Hex Addr	1720	5920
x"00",	-- Hex Addr	1721	5921
x"00",	-- Hex Addr	1722	5922
x"00",	-- Hex Addr	1723	5923
x"00",	-- Hex Addr	1724	5924
x"00",	-- Hex Addr	1725	5925
x"00",	-- Hex Addr	1726	5926
x"00",	-- Hex Addr	1727	5927
x"00",	-- Hex Addr	1728	5928
x"00",	-- Hex Addr	1729	5929
x"00",	-- Hex Addr	172A	5930
x"00",	-- Hex Addr	172B	5931
x"00",	-- Hex Addr	172C	5932
x"00",	-- Hex Addr	172D	5933
x"00",	-- Hex Addr	172E	5934
x"00",	-- Hex Addr	172F	5935
x"00",	-- Hex Addr	1730	5936
x"00",	-- Hex Addr	1731	5937
x"00",	-- Hex Addr	1732	5938
x"00",	-- Hex Addr	1733	5939
x"00",	-- Hex Addr	1734	5940
x"00",	-- Hex Addr	1735	5941
x"00",	-- Hex Addr	1736	5942
x"00",	-- Hex Addr	1737	5943
x"00",	-- Hex Addr	1738	5944
x"00",	-- Hex Addr	1739	5945
x"00",	-- Hex Addr	173A	5946
x"00",	-- Hex Addr	173B	5947
x"00",	-- Hex Addr	173C	5948
x"00",	-- Hex Addr	173D	5949
x"00",	-- Hex Addr	173E	5950
x"00",	-- Hex Addr	173F	5951
x"00",	-- Hex Addr	1740	5952
x"00",	-- Hex Addr	1741	5953
x"00",	-- Hex Addr	1742	5954
x"00",	-- Hex Addr	1743	5955
x"00",	-- Hex Addr	1744	5956
x"00",	-- Hex Addr	1745	5957
x"00",	-- Hex Addr	1746	5958
x"00",	-- Hex Addr	1747	5959
x"00",	-- Hex Addr	1748	5960
x"00",	-- Hex Addr	1749	5961
x"00",	-- Hex Addr	174A	5962
x"00",	-- Hex Addr	174B	5963
x"00",	-- Hex Addr	174C	5964
x"00",	-- Hex Addr	174D	5965
x"00",	-- Hex Addr	174E	5966
x"00",	-- Hex Addr	174F	5967
x"00",	-- Hex Addr	1750	5968
x"00",	-- Hex Addr	1751	5969
x"00",	-- Hex Addr	1752	5970
x"00",	-- Hex Addr	1753	5971
x"00",	-- Hex Addr	1754	5972
x"00",	-- Hex Addr	1755	5973
x"00",	-- Hex Addr	1756	5974
x"00",	-- Hex Addr	1757	5975
x"00",	-- Hex Addr	1758	5976
x"00",	-- Hex Addr	1759	5977
x"00",	-- Hex Addr	175A	5978
x"00",	-- Hex Addr	175B	5979
x"00",	-- Hex Addr	175C	5980
x"00",	-- Hex Addr	175D	5981
x"00",	-- Hex Addr	175E	5982
x"00",	-- Hex Addr	175F	5983
x"00",	-- Hex Addr	1760	5984
x"00",	-- Hex Addr	1761	5985
x"00",	-- Hex Addr	1762	5986
x"00",	-- Hex Addr	1763	5987
x"00",	-- Hex Addr	1764	5988
x"00",	-- Hex Addr	1765	5989
x"00",	-- Hex Addr	1766	5990
x"00",	-- Hex Addr	1767	5991
x"00",	-- Hex Addr	1768	5992
x"00",	-- Hex Addr	1769	5993
x"00",	-- Hex Addr	176A	5994
x"00",	-- Hex Addr	176B	5995
x"00",	-- Hex Addr	176C	5996
x"00",	-- Hex Addr	176D	5997
x"00",	-- Hex Addr	176E	5998
x"00",	-- Hex Addr	176F	5999
x"00",	-- Hex Addr	1770	6000
x"00",	-- Hex Addr	1771	6001
x"00",	-- Hex Addr	1772	6002
x"00",	-- Hex Addr	1773	6003
x"00",	-- Hex Addr	1774	6004
x"00",	-- Hex Addr	1775	6005
x"00",	-- Hex Addr	1776	6006
x"00",	-- Hex Addr	1777	6007
x"00",	-- Hex Addr	1778	6008
x"00",	-- Hex Addr	1779	6009
x"00",	-- Hex Addr	177A	6010
x"00",	-- Hex Addr	177B	6011
x"00",	-- Hex Addr	177C	6012
x"00",	-- Hex Addr	177D	6013
x"00",	-- Hex Addr	177E	6014
x"00",	-- Hex Addr	177F	6015
x"00",	-- Hex Addr	1780	6016
x"00",	-- Hex Addr	1781	6017
x"00",	-- Hex Addr	1782	6018
x"00",	-- Hex Addr	1783	6019
x"00",	-- Hex Addr	1784	6020
x"00",	-- Hex Addr	1785	6021
x"00",	-- Hex Addr	1786	6022
x"00",	-- Hex Addr	1787	6023
x"00",	-- Hex Addr	1788	6024
x"00",	-- Hex Addr	1789	6025
x"00",	-- Hex Addr	178A	6026
x"00",	-- Hex Addr	178B	6027
x"00",	-- Hex Addr	178C	6028
x"00",	-- Hex Addr	178D	6029
x"00",	-- Hex Addr	178E	6030
x"00",	-- Hex Addr	178F	6031
x"00",	-- Hex Addr	1790	6032
x"00",	-- Hex Addr	1791	6033
x"00",	-- Hex Addr	1792	6034
x"00",	-- Hex Addr	1793	6035
x"00",	-- Hex Addr	1794	6036
x"00",	-- Hex Addr	1795	6037
x"00",	-- Hex Addr	1796	6038
x"00",	-- Hex Addr	1797	6039
x"00",	-- Hex Addr	1798	6040
x"00",	-- Hex Addr	1799	6041
x"00",	-- Hex Addr	179A	6042
x"00",	-- Hex Addr	179B	6043
x"00",	-- Hex Addr	179C	6044
x"00",	-- Hex Addr	179D	6045
x"00",	-- Hex Addr	179E	6046
x"00",	-- Hex Addr	179F	6047
x"00",	-- Hex Addr	17A0	6048
x"00",	-- Hex Addr	17A1	6049
x"00",	-- Hex Addr	17A2	6050
x"00",	-- Hex Addr	17A3	6051
x"00",	-- Hex Addr	17A4	6052
x"00",	-- Hex Addr	17A5	6053
x"00",	-- Hex Addr	17A6	6054
x"00",	-- Hex Addr	17A7	6055
x"00",	-- Hex Addr	17A8	6056
x"00",	-- Hex Addr	17A9	6057
x"00",	-- Hex Addr	17AA	6058
x"00",	-- Hex Addr	17AB	6059
x"00",	-- Hex Addr	17AC	6060
x"00",	-- Hex Addr	17AD	6061
x"00",	-- Hex Addr	17AE	6062
x"00",	-- Hex Addr	17AF	6063
x"00",	-- Hex Addr	17B0	6064
x"00",	-- Hex Addr	17B1	6065
x"00",	-- Hex Addr	17B2	6066
x"00",	-- Hex Addr	17B3	6067
x"00",	-- Hex Addr	17B4	6068
x"00",	-- Hex Addr	17B5	6069
x"00",	-- Hex Addr	17B6	6070
x"00",	-- Hex Addr	17B7	6071
x"00",	-- Hex Addr	17B8	6072
x"00",	-- Hex Addr	17B9	6073
x"00",	-- Hex Addr	17BA	6074
x"00",	-- Hex Addr	17BB	6075
x"00",	-- Hex Addr	17BC	6076
x"00",	-- Hex Addr	17BD	6077
x"00",	-- Hex Addr	17BE	6078
x"00",	-- Hex Addr	17BF	6079
x"00",	-- Hex Addr	17C0	6080
x"00",	-- Hex Addr	17C1	6081
x"00",	-- Hex Addr	17C2	6082
x"00",	-- Hex Addr	17C3	6083
x"00",	-- Hex Addr	17C4	6084
x"00",	-- Hex Addr	17C5	6085
x"00",	-- Hex Addr	17C6	6086
x"00",	-- Hex Addr	17C7	6087
x"00",	-- Hex Addr	17C8	6088
x"00",	-- Hex Addr	17C9	6089
x"00",	-- Hex Addr	17CA	6090
x"00",	-- Hex Addr	17CB	6091
x"00",	-- Hex Addr	17CC	6092
x"00",	-- Hex Addr	17CD	6093
x"00",	-- Hex Addr	17CE	6094
x"00",	-- Hex Addr	17CF	6095
x"00",	-- Hex Addr	17D0	6096
x"00",	-- Hex Addr	17D1	6097
x"00",	-- Hex Addr	17D2	6098
x"00",	-- Hex Addr	17D3	6099
x"00",	-- Hex Addr	17D4	6100
x"00",	-- Hex Addr	17D5	6101
x"00",	-- Hex Addr	17D6	6102
x"00",	-- Hex Addr	17D7	6103
x"00",	-- Hex Addr	17D8	6104
x"00",	-- Hex Addr	17D9	6105
x"00",	-- Hex Addr	17DA	6106
x"00",	-- Hex Addr	17DB	6107
x"00",	-- Hex Addr	17DC	6108
x"00",	-- Hex Addr	17DD	6109
x"00",	-- Hex Addr	17DE	6110
x"00",	-- Hex Addr	17DF	6111
x"00",	-- Hex Addr	17E0	6112
x"00",	-- Hex Addr	17E1	6113
x"00",	-- Hex Addr	17E2	6114
x"00",	-- Hex Addr	17E3	6115
x"00",	-- Hex Addr	17E4	6116
x"00",	-- Hex Addr	17E5	6117
x"00",	-- Hex Addr	17E6	6118
x"00",	-- Hex Addr	17E7	6119
x"00",	-- Hex Addr	17E8	6120
x"00",	-- Hex Addr	17E9	6121
x"00",	-- Hex Addr	17EA	6122
x"00",	-- Hex Addr	17EB	6123
x"00",	-- Hex Addr	17EC	6124
x"00",	-- Hex Addr	17ED	6125
x"00",	-- Hex Addr	17EE	6126
x"00",	-- Hex Addr	17EF	6127
x"00",	-- Hex Addr	17F0	6128
x"00",	-- Hex Addr	17F1	6129
x"00",	-- Hex Addr	17F2	6130
x"00",	-- Hex Addr	17F3	6131
x"00",	-- Hex Addr	17F4	6132
x"00",	-- Hex Addr	17F5	6133
x"00",	-- Hex Addr	17F6	6134
x"00",	-- Hex Addr	17F7	6135
x"00",	-- Hex Addr	17F8	6136
x"00",	-- Hex Addr	17F9	6137
x"00",	-- Hex Addr	17FA	6138
x"00",	-- Hex Addr	17FB	6139
x"00",	-- Hex Addr	17FC	6140
x"00",	-- Hex Addr	17FD	6141
x"00",	-- Hex Addr	17FE	6142
x"00",	-- Hex Addr	17FF	6143
x"00",	-- Hex Addr	1800	6144
x"00",	-- Hex Addr	1801	6145
x"00",	-- Hex Addr	1802	6146
x"00",	-- Hex Addr	1803	6147
x"00",	-- Hex Addr	1804	6148
x"00",	-- Hex Addr	1805	6149
x"00",	-- Hex Addr	1806	6150
x"00",	-- Hex Addr	1807	6151
x"00",	-- Hex Addr	1808	6152
x"00",	-- Hex Addr	1809	6153
x"00",	-- Hex Addr	180A	6154
x"00",	-- Hex Addr	180B	6155
x"00",	-- Hex Addr	180C	6156
x"00",	-- Hex Addr	180D	6157
x"00",	-- Hex Addr	180E	6158
x"00",	-- Hex Addr	180F	6159
x"00",	-- Hex Addr	1810	6160
x"00",	-- Hex Addr	1811	6161
x"00",	-- Hex Addr	1812	6162
x"00",	-- Hex Addr	1813	6163
x"00",	-- Hex Addr	1814	6164
x"00",	-- Hex Addr	1815	6165
x"00",	-- Hex Addr	1816	6166
x"00",	-- Hex Addr	1817	6167
x"00",	-- Hex Addr	1818	6168
x"00",	-- Hex Addr	1819	6169
x"00",	-- Hex Addr	181A	6170
x"00",	-- Hex Addr	181B	6171
x"00",	-- Hex Addr	181C	6172
x"00",	-- Hex Addr	181D	6173
x"00",	-- Hex Addr	181E	6174
x"00",	-- Hex Addr	181F	6175
x"00",	-- Hex Addr	1820	6176
x"00",	-- Hex Addr	1821	6177
x"00",	-- Hex Addr	1822	6178
x"00",	-- Hex Addr	1823	6179
x"00",	-- Hex Addr	1824	6180
x"00",	-- Hex Addr	1825	6181
x"00",	-- Hex Addr	1826	6182
x"00",	-- Hex Addr	1827	6183
x"00",	-- Hex Addr	1828	6184
x"00",	-- Hex Addr	1829	6185
x"00",	-- Hex Addr	182A	6186
x"00",	-- Hex Addr	182B	6187
x"00",	-- Hex Addr	182C	6188
x"00",	-- Hex Addr	182D	6189
x"00",	-- Hex Addr	182E	6190
x"00",	-- Hex Addr	182F	6191
x"00",	-- Hex Addr	1830	6192
x"00",	-- Hex Addr	1831	6193
x"00",	-- Hex Addr	1832	6194
x"00",	-- Hex Addr	1833	6195
x"00",	-- Hex Addr	1834	6196
x"00",	-- Hex Addr	1835	6197
x"00",	-- Hex Addr	1836	6198
x"00",	-- Hex Addr	1837	6199
x"00",	-- Hex Addr	1838	6200
x"00",	-- Hex Addr	1839	6201
x"00",	-- Hex Addr	183A	6202
x"00",	-- Hex Addr	183B	6203
x"00",	-- Hex Addr	183C	6204
x"00",	-- Hex Addr	183D	6205
x"00",	-- Hex Addr	183E	6206
x"00",	-- Hex Addr	183F	6207
x"00",	-- Hex Addr	1840	6208
x"00",	-- Hex Addr	1841	6209
x"00",	-- Hex Addr	1842	6210
x"00",	-- Hex Addr	1843	6211
x"00",	-- Hex Addr	1844	6212
x"00",	-- Hex Addr	1845	6213
x"00",	-- Hex Addr	1846	6214
x"00",	-- Hex Addr	1847	6215
x"00",	-- Hex Addr	1848	6216
x"00",	-- Hex Addr	1849	6217
x"00",	-- Hex Addr	184A	6218
x"00",	-- Hex Addr	184B	6219
x"00",	-- Hex Addr	184C	6220
x"00",	-- Hex Addr	184D	6221
x"00",	-- Hex Addr	184E	6222
x"00",	-- Hex Addr	184F	6223
x"00",	-- Hex Addr	1850	6224
x"00",	-- Hex Addr	1851	6225
x"00",	-- Hex Addr	1852	6226
x"00",	-- Hex Addr	1853	6227
x"00",	-- Hex Addr	1854	6228
x"00",	-- Hex Addr	1855	6229
x"00",	-- Hex Addr	1856	6230
x"00",	-- Hex Addr	1857	6231
x"00",	-- Hex Addr	1858	6232
x"00",	-- Hex Addr	1859	6233
x"00",	-- Hex Addr	185A	6234
x"00",	-- Hex Addr	185B	6235
x"00",	-- Hex Addr	185C	6236
x"00",	-- Hex Addr	185D	6237
x"00",	-- Hex Addr	185E	6238
x"00",	-- Hex Addr	185F	6239
x"00",	-- Hex Addr	1860	6240
x"00",	-- Hex Addr	1861	6241
x"00",	-- Hex Addr	1862	6242
x"00",	-- Hex Addr	1863	6243
x"00",	-- Hex Addr	1864	6244
x"00",	-- Hex Addr	1865	6245
x"00",	-- Hex Addr	1866	6246
x"00",	-- Hex Addr	1867	6247
x"00",	-- Hex Addr	1868	6248
x"00",	-- Hex Addr	1869	6249
x"00",	-- Hex Addr	186A	6250
x"00",	-- Hex Addr	186B	6251
x"00",	-- Hex Addr	186C	6252
x"00",	-- Hex Addr	186D	6253
x"00",	-- Hex Addr	186E	6254
x"00",	-- Hex Addr	186F	6255
x"00",	-- Hex Addr	1870	6256
x"00",	-- Hex Addr	1871	6257
x"00",	-- Hex Addr	1872	6258
x"00",	-- Hex Addr	1873	6259
x"00",	-- Hex Addr	1874	6260
x"00",	-- Hex Addr	1875	6261
x"00",	-- Hex Addr	1876	6262
x"00",	-- Hex Addr	1877	6263
x"00",	-- Hex Addr	1878	6264
x"00",	-- Hex Addr	1879	6265
x"00",	-- Hex Addr	187A	6266
x"00",	-- Hex Addr	187B	6267
x"00",	-- Hex Addr	187C	6268
x"00",	-- Hex Addr	187D	6269
x"00",	-- Hex Addr	187E	6270
x"00",	-- Hex Addr	187F	6271
x"00",	-- Hex Addr	1880	6272
x"00",	-- Hex Addr	1881	6273
x"00",	-- Hex Addr	1882	6274
x"00",	-- Hex Addr	1883	6275
x"00",	-- Hex Addr	1884	6276
x"00",	-- Hex Addr	1885	6277
x"00",	-- Hex Addr	1886	6278
x"00",	-- Hex Addr	1887	6279
x"00",	-- Hex Addr	1888	6280
x"00",	-- Hex Addr	1889	6281
x"00",	-- Hex Addr	188A	6282
x"00",	-- Hex Addr	188B	6283
x"00",	-- Hex Addr	188C	6284
x"00",	-- Hex Addr	188D	6285
x"00",	-- Hex Addr	188E	6286
x"00",	-- Hex Addr	188F	6287
x"00",	-- Hex Addr	1890	6288
x"00",	-- Hex Addr	1891	6289
x"00",	-- Hex Addr	1892	6290
x"00",	-- Hex Addr	1893	6291
x"00",	-- Hex Addr	1894	6292
x"00",	-- Hex Addr	1895	6293
x"00",	-- Hex Addr	1896	6294
x"00",	-- Hex Addr	1897	6295
x"00",	-- Hex Addr	1898	6296
x"00",	-- Hex Addr	1899	6297
x"00",	-- Hex Addr	189A	6298
x"00",	-- Hex Addr	189B	6299
x"00",	-- Hex Addr	189C	6300
x"00",	-- Hex Addr	189D	6301
x"00",	-- Hex Addr	189E	6302
x"00",	-- Hex Addr	189F	6303
x"00",	-- Hex Addr	18A0	6304
x"00",	-- Hex Addr	18A1	6305
x"00",	-- Hex Addr	18A2	6306
x"00",	-- Hex Addr	18A3	6307
x"00",	-- Hex Addr	18A4	6308
x"00",	-- Hex Addr	18A5	6309
x"00",	-- Hex Addr	18A6	6310
x"00",	-- Hex Addr	18A7	6311
x"00",	-- Hex Addr	18A8	6312
x"00",	-- Hex Addr	18A9	6313
x"00",	-- Hex Addr	18AA	6314
x"00",	-- Hex Addr	18AB	6315
x"00",	-- Hex Addr	18AC	6316
x"00",	-- Hex Addr	18AD	6317
x"00",	-- Hex Addr	18AE	6318
x"00",	-- Hex Addr	18AF	6319
x"00",	-- Hex Addr	18B0	6320
x"00",	-- Hex Addr	18B1	6321
x"00",	-- Hex Addr	18B2	6322
x"00",	-- Hex Addr	18B3	6323
x"00",	-- Hex Addr	18B4	6324
x"00",	-- Hex Addr	18B5	6325
x"00",	-- Hex Addr	18B6	6326
x"00",	-- Hex Addr	18B7	6327
x"00",	-- Hex Addr	18B8	6328
x"00",	-- Hex Addr	18B9	6329
x"00",	-- Hex Addr	18BA	6330
x"00",	-- Hex Addr	18BB	6331
x"00",	-- Hex Addr	18BC	6332
x"00",	-- Hex Addr	18BD	6333
x"00",	-- Hex Addr	18BE	6334
x"00",	-- Hex Addr	18BF	6335
x"00",	-- Hex Addr	18C0	6336
x"00",	-- Hex Addr	18C1	6337
x"00",	-- Hex Addr	18C2	6338
x"00",	-- Hex Addr	18C3	6339
x"00",	-- Hex Addr	18C4	6340
x"00",	-- Hex Addr	18C5	6341
x"00",	-- Hex Addr	18C6	6342
x"00",	-- Hex Addr	18C7	6343
x"00",	-- Hex Addr	18C8	6344
x"00",	-- Hex Addr	18C9	6345
x"00",	-- Hex Addr	18CA	6346
x"00",	-- Hex Addr	18CB	6347
x"00",	-- Hex Addr	18CC	6348
x"00",	-- Hex Addr	18CD	6349
x"00",	-- Hex Addr	18CE	6350
x"00",	-- Hex Addr	18CF	6351
x"00",	-- Hex Addr	18D0	6352
x"00",	-- Hex Addr	18D1	6353
x"00",	-- Hex Addr	18D2	6354
x"00",	-- Hex Addr	18D3	6355
x"00",	-- Hex Addr	18D4	6356
x"00",	-- Hex Addr	18D5	6357
x"00",	-- Hex Addr	18D6	6358
x"00",	-- Hex Addr	18D7	6359
x"00",	-- Hex Addr	18D8	6360
x"00",	-- Hex Addr	18D9	6361
x"00",	-- Hex Addr	18DA	6362
x"00",	-- Hex Addr	18DB	6363
x"00",	-- Hex Addr	18DC	6364
x"00",	-- Hex Addr	18DD	6365
x"00",	-- Hex Addr	18DE	6366
x"00",	-- Hex Addr	18DF	6367
x"00",	-- Hex Addr	18E0	6368
x"00",	-- Hex Addr	18E1	6369
x"00",	-- Hex Addr	18E2	6370
x"00",	-- Hex Addr	18E3	6371
x"00",	-- Hex Addr	18E4	6372
x"00",	-- Hex Addr	18E5	6373
x"00",	-- Hex Addr	18E6	6374
x"00",	-- Hex Addr	18E7	6375
x"00",	-- Hex Addr	18E8	6376
x"00",	-- Hex Addr	18E9	6377
x"00",	-- Hex Addr	18EA	6378
x"00",	-- Hex Addr	18EB	6379
x"00",	-- Hex Addr	18EC	6380
x"00",	-- Hex Addr	18ED	6381
x"00",	-- Hex Addr	18EE	6382
x"00",	-- Hex Addr	18EF	6383
x"00",	-- Hex Addr	18F0	6384
x"00",	-- Hex Addr	18F1	6385
x"00",	-- Hex Addr	18F2	6386
x"00",	-- Hex Addr	18F3	6387
x"00",	-- Hex Addr	18F4	6388
x"00",	-- Hex Addr	18F5	6389
x"00",	-- Hex Addr	18F6	6390
x"00",	-- Hex Addr	18F7	6391
x"00",	-- Hex Addr	18F8	6392
x"00",	-- Hex Addr	18F9	6393
x"00",	-- Hex Addr	18FA	6394
x"00",	-- Hex Addr	18FB	6395
x"00",	-- Hex Addr	18FC	6396
x"00",	-- Hex Addr	18FD	6397
x"00",	-- Hex Addr	18FE	6398
x"00",	-- Hex Addr	18FF	6399
x"00",	-- Hex Addr	1900	6400
x"00",	-- Hex Addr	1901	6401
x"00",	-- Hex Addr	1902	6402
x"00",	-- Hex Addr	1903	6403
x"00",	-- Hex Addr	1904	6404
x"00",	-- Hex Addr	1905	6405
x"00",	-- Hex Addr	1906	6406
x"00",	-- Hex Addr	1907	6407
x"00",	-- Hex Addr	1908	6408
x"00",	-- Hex Addr	1909	6409
x"00",	-- Hex Addr	190A	6410
x"00",	-- Hex Addr	190B	6411
x"00",	-- Hex Addr	190C	6412
x"00",	-- Hex Addr	190D	6413
x"00",	-- Hex Addr	190E	6414
x"00",	-- Hex Addr	190F	6415
x"00",	-- Hex Addr	1910	6416
x"00",	-- Hex Addr	1911	6417
x"00",	-- Hex Addr	1912	6418
x"00",	-- Hex Addr	1913	6419
x"00",	-- Hex Addr	1914	6420
x"00",	-- Hex Addr	1915	6421
x"00",	-- Hex Addr	1916	6422
x"00",	-- Hex Addr	1917	6423
x"00",	-- Hex Addr	1918	6424
x"00",	-- Hex Addr	1919	6425
x"00",	-- Hex Addr	191A	6426
x"00",	-- Hex Addr	191B	6427
x"00",	-- Hex Addr	191C	6428
x"00",	-- Hex Addr	191D	6429
x"00",	-- Hex Addr	191E	6430
x"00",	-- Hex Addr	191F	6431
x"00",	-- Hex Addr	1920	6432
x"00",	-- Hex Addr	1921	6433
x"00",	-- Hex Addr	1922	6434
x"00",	-- Hex Addr	1923	6435
x"00",	-- Hex Addr	1924	6436
x"00",	-- Hex Addr	1925	6437
x"00",	-- Hex Addr	1926	6438
x"00",	-- Hex Addr	1927	6439
x"00",	-- Hex Addr	1928	6440
x"00",	-- Hex Addr	1929	6441
x"00",	-- Hex Addr	192A	6442
x"00",	-- Hex Addr	192B	6443
x"00",	-- Hex Addr	192C	6444
x"00",	-- Hex Addr	192D	6445
x"00",	-- Hex Addr	192E	6446
x"00",	-- Hex Addr	192F	6447
x"00",	-- Hex Addr	1930	6448
x"00",	-- Hex Addr	1931	6449
x"00",	-- Hex Addr	1932	6450
x"00",	-- Hex Addr	1933	6451
x"00",	-- Hex Addr	1934	6452
x"00",	-- Hex Addr	1935	6453
x"00",	-- Hex Addr	1936	6454
x"00",	-- Hex Addr	1937	6455
x"00",	-- Hex Addr	1938	6456
x"00",	-- Hex Addr	1939	6457
x"00",	-- Hex Addr	193A	6458
x"00",	-- Hex Addr	193B	6459
x"00",	-- Hex Addr	193C	6460
x"00",	-- Hex Addr	193D	6461
x"00",	-- Hex Addr	193E	6462
x"00",	-- Hex Addr	193F	6463
x"00",	-- Hex Addr	1940	6464
x"00",	-- Hex Addr	1941	6465
x"00",	-- Hex Addr	1942	6466
x"00",	-- Hex Addr	1943	6467
x"00",	-- Hex Addr	1944	6468
x"00",	-- Hex Addr	1945	6469
x"00",	-- Hex Addr	1946	6470
x"00",	-- Hex Addr	1947	6471
x"00",	-- Hex Addr	1948	6472
x"00",	-- Hex Addr	1949	6473
x"00",	-- Hex Addr	194A	6474
x"00",	-- Hex Addr	194B	6475
x"00",	-- Hex Addr	194C	6476
x"00",	-- Hex Addr	194D	6477
x"00",	-- Hex Addr	194E	6478
x"00",	-- Hex Addr	194F	6479
x"00",	-- Hex Addr	1950	6480
x"00",	-- Hex Addr	1951	6481
x"00",	-- Hex Addr	1952	6482
x"00",	-- Hex Addr	1953	6483
x"00",	-- Hex Addr	1954	6484
x"00",	-- Hex Addr	1955	6485
x"00",	-- Hex Addr	1956	6486
x"00",	-- Hex Addr	1957	6487
x"00",	-- Hex Addr	1958	6488
x"00",	-- Hex Addr	1959	6489
x"00",	-- Hex Addr	195A	6490
x"00",	-- Hex Addr	195B	6491
x"00",	-- Hex Addr	195C	6492
x"00",	-- Hex Addr	195D	6493
x"00",	-- Hex Addr	195E	6494
x"00",	-- Hex Addr	195F	6495
x"00",	-- Hex Addr	1960	6496
x"00",	-- Hex Addr	1961	6497
x"00",	-- Hex Addr	1962	6498
x"00",	-- Hex Addr	1963	6499
x"00",	-- Hex Addr	1964	6500
x"00",	-- Hex Addr	1965	6501
x"00",	-- Hex Addr	1966	6502
x"00",	-- Hex Addr	1967	6503
x"00",	-- Hex Addr	1968	6504
x"00",	-- Hex Addr	1969	6505
x"00",	-- Hex Addr	196A	6506
x"00",	-- Hex Addr	196B	6507
x"00",	-- Hex Addr	196C	6508
x"00",	-- Hex Addr	196D	6509
x"00",	-- Hex Addr	196E	6510
x"00",	-- Hex Addr	196F	6511
x"00",	-- Hex Addr	1970	6512
x"00",	-- Hex Addr	1971	6513
x"00",	-- Hex Addr	1972	6514
x"00",	-- Hex Addr	1973	6515
x"00",	-- Hex Addr	1974	6516
x"00",	-- Hex Addr	1975	6517
x"00",	-- Hex Addr	1976	6518
x"00",	-- Hex Addr	1977	6519
x"00",	-- Hex Addr	1978	6520
x"00",	-- Hex Addr	1979	6521
x"00",	-- Hex Addr	197A	6522
x"00",	-- Hex Addr	197B	6523
x"00",	-- Hex Addr	197C	6524
x"00",	-- Hex Addr	197D	6525
x"00",	-- Hex Addr	197E	6526
x"00",	-- Hex Addr	197F	6527
x"00",	-- Hex Addr	1980	6528
x"00",	-- Hex Addr	1981	6529
x"00",	-- Hex Addr	1982	6530
x"00",	-- Hex Addr	1983	6531
x"00",	-- Hex Addr	1984	6532
x"00",	-- Hex Addr	1985	6533
x"00",	-- Hex Addr	1986	6534
x"00",	-- Hex Addr	1987	6535
x"00",	-- Hex Addr	1988	6536
x"00",	-- Hex Addr	1989	6537
x"00",	-- Hex Addr	198A	6538
x"00",	-- Hex Addr	198B	6539
x"00",	-- Hex Addr	198C	6540
x"00",	-- Hex Addr	198D	6541
x"00",	-- Hex Addr	198E	6542
x"00",	-- Hex Addr	198F	6543
x"00",	-- Hex Addr	1990	6544
x"00",	-- Hex Addr	1991	6545
x"00",	-- Hex Addr	1992	6546
x"00",	-- Hex Addr	1993	6547
x"00",	-- Hex Addr	1994	6548
x"00",	-- Hex Addr	1995	6549
x"00",	-- Hex Addr	1996	6550
x"00",	-- Hex Addr	1997	6551
x"00",	-- Hex Addr	1998	6552
x"00",	-- Hex Addr	1999	6553
x"00",	-- Hex Addr	199A	6554
x"00",	-- Hex Addr	199B	6555
x"00",	-- Hex Addr	199C	6556
x"00",	-- Hex Addr	199D	6557
x"00",	-- Hex Addr	199E	6558
x"00",	-- Hex Addr	199F	6559
x"00",	-- Hex Addr	19A0	6560
x"00",	-- Hex Addr	19A1	6561
x"00",	-- Hex Addr	19A2	6562
x"00",	-- Hex Addr	19A3	6563
x"00",	-- Hex Addr	19A4	6564
x"00",	-- Hex Addr	19A5	6565
x"00",	-- Hex Addr	19A6	6566
x"00",	-- Hex Addr	19A7	6567
x"00",	-- Hex Addr	19A8	6568
x"00",	-- Hex Addr	19A9	6569
x"00",	-- Hex Addr	19AA	6570
x"00",	-- Hex Addr	19AB	6571
x"00",	-- Hex Addr	19AC	6572
x"00",	-- Hex Addr	19AD	6573
x"00",	-- Hex Addr	19AE	6574
x"00",	-- Hex Addr	19AF	6575
x"00",	-- Hex Addr	19B0	6576
x"00",	-- Hex Addr	19B1	6577
x"00",	-- Hex Addr	19B2	6578
x"00",	-- Hex Addr	19B3	6579
x"00",	-- Hex Addr	19B4	6580
x"00",	-- Hex Addr	19B5	6581
x"00",	-- Hex Addr	19B6	6582
x"00",	-- Hex Addr	19B7	6583
x"00",	-- Hex Addr	19B8	6584
x"00",	-- Hex Addr	19B9	6585
x"00",	-- Hex Addr	19BA	6586
x"00",	-- Hex Addr	19BB	6587
x"00",	-- Hex Addr	19BC	6588
x"00",	-- Hex Addr	19BD	6589
x"00",	-- Hex Addr	19BE	6590
x"00",	-- Hex Addr	19BF	6591
x"00",	-- Hex Addr	19C0	6592
x"00",	-- Hex Addr	19C1	6593
x"00",	-- Hex Addr	19C2	6594
x"00",	-- Hex Addr	19C3	6595
x"00",	-- Hex Addr	19C4	6596
x"00",	-- Hex Addr	19C5	6597
x"00",	-- Hex Addr	19C6	6598
x"00",	-- Hex Addr	19C7	6599
x"00",	-- Hex Addr	19C8	6600
x"00",	-- Hex Addr	19C9	6601
x"00",	-- Hex Addr	19CA	6602
x"00",	-- Hex Addr	19CB	6603
x"00",	-- Hex Addr	19CC	6604
x"00",	-- Hex Addr	19CD	6605
x"00",	-- Hex Addr	19CE	6606
x"00",	-- Hex Addr	19CF	6607
x"00",	-- Hex Addr	19D0	6608
x"00",	-- Hex Addr	19D1	6609
x"00",	-- Hex Addr	19D2	6610
x"00",	-- Hex Addr	19D3	6611
x"00",	-- Hex Addr	19D4	6612
x"00",	-- Hex Addr	19D5	6613
x"00",	-- Hex Addr	19D6	6614
x"00",	-- Hex Addr	19D7	6615
x"00",	-- Hex Addr	19D8	6616
x"00",	-- Hex Addr	19D9	6617
x"00",	-- Hex Addr	19DA	6618
x"00",	-- Hex Addr	19DB	6619
x"00",	-- Hex Addr	19DC	6620
x"00",	-- Hex Addr	19DD	6621
x"00",	-- Hex Addr	19DE	6622
x"00",	-- Hex Addr	19DF	6623
x"00",	-- Hex Addr	19E0	6624
x"00",	-- Hex Addr	19E1	6625
x"00",	-- Hex Addr	19E2	6626
x"00",	-- Hex Addr	19E3	6627
x"00",	-- Hex Addr	19E4	6628
x"00",	-- Hex Addr	19E5	6629
x"00",	-- Hex Addr	19E6	6630
x"00",	-- Hex Addr	19E7	6631
x"00",	-- Hex Addr	19E8	6632
x"00",	-- Hex Addr	19E9	6633
x"00",	-- Hex Addr	19EA	6634
x"00",	-- Hex Addr	19EB	6635
x"00",	-- Hex Addr	19EC	6636
x"00",	-- Hex Addr	19ED	6637
x"00",	-- Hex Addr	19EE	6638
x"00",	-- Hex Addr	19EF	6639
x"00",	-- Hex Addr	19F0	6640
x"00",	-- Hex Addr	19F1	6641
x"00",	-- Hex Addr	19F2	6642
x"00",	-- Hex Addr	19F3	6643
x"00",	-- Hex Addr	19F4	6644
x"00",	-- Hex Addr	19F5	6645
x"00",	-- Hex Addr	19F6	6646
x"00",	-- Hex Addr	19F7	6647
x"00",	-- Hex Addr	19F8	6648
x"00",	-- Hex Addr	19F9	6649
x"00",	-- Hex Addr	19FA	6650
x"00",	-- Hex Addr	19FB	6651
x"00",	-- Hex Addr	19FC	6652
x"00",	-- Hex Addr	19FD	6653
x"00",	-- Hex Addr	19FE	6654
x"00",	-- Hex Addr	19FF	6655
x"00",	-- Hex Addr	1A00	6656
x"00",	-- Hex Addr	1A01	6657
x"00",	-- Hex Addr	1A02	6658
x"00",	-- Hex Addr	1A03	6659
x"00",	-- Hex Addr	1A04	6660
x"00",	-- Hex Addr	1A05	6661
x"00",	-- Hex Addr	1A06	6662
x"00",	-- Hex Addr	1A07	6663
x"00",	-- Hex Addr	1A08	6664
x"00",	-- Hex Addr	1A09	6665
x"00",	-- Hex Addr	1A0A	6666
x"00",	-- Hex Addr	1A0B	6667
x"00",	-- Hex Addr	1A0C	6668
x"00",	-- Hex Addr	1A0D	6669
x"00",	-- Hex Addr	1A0E	6670
x"00",	-- Hex Addr	1A0F	6671
x"00",	-- Hex Addr	1A10	6672
x"00",	-- Hex Addr	1A11	6673
x"00",	-- Hex Addr	1A12	6674
x"00",	-- Hex Addr	1A13	6675
x"00",	-- Hex Addr	1A14	6676
x"00",	-- Hex Addr	1A15	6677
x"00",	-- Hex Addr	1A16	6678
x"00",	-- Hex Addr	1A17	6679
x"00",	-- Hex Addr	1A18	6680
x"00",	-- Hex Addr	1A19	6681
x"00",	-- Hex Addr	1A1A	6682
x"00",	-- Hex Addr	1A1B	6683
x"00",	-- Hex Addr	1A1C	6684
x"00",	-- Hex Addr	1A1D	6685
x"00",	-- Hex Addr	1A1E	6686
x"00",	-- Hex Addr	1A1F	6687
x"00",	-- Hex Addr	1A20	6688
x"00",	-- Hex Addr	1A21	6689
x"00",	-- Hex Addr	1A22	6690
x"00",	-- Hex Addr	1A23	6691
x"00",	-- Hex Addr	1A24	6692
x"00",	-- Hex Addr	1A25	6693
x"00",	-- Hex Addr	1A26	6694
x"00",	-- Hex Addr	1A27	6695
x"00",	-- Hex Addr	1A28	6696
x"00",	-- Hex Addr	1A29	6697
x"00",	-- Hex Addr	1A2A	6698
x"00",	-- Hex Addr	1A2B	6699
x"00",	-- Hex Addr	1A2C	6700
x"00",	-- Hex Addr	1A2D	6701
x"00",	-- Hex Addr	1A2E	6702
x"00",	-- Hex Addr	1A2F	6703
x"00",	-- Hex Addr	1A30	6704
x"00",	-- Hex Addr	1A31	6705
x"00",	-- Hex Addr	1A32	6706
x"00",	-- Hex Addr	1A33	6707
x"00",	-- Hex Addr	1A34	6708
x"00",	-- Hex Addr	1A35	6709
x"00",	-- Hex Addr	1A36	6710
x"00",	-- Hex Addr	1A37	6711
x"00",	-- Hex Addr	1A38	6712
x"00",	-- Hex Addr	1A39	6713
x"00",	-- Hex Addr	1A3A	6714
x"00",	-- Hex Addr	1A3B	6715
x"00",	-- Hex Addr	1A3C	6716
x"00",	-- Hex Addr	1A3D	6717
x"00",	-- Hex Addr	1A3E	6718
x"00",	-- Hex Addr	1A3F	6719
x"00",	-- Hex Addr	1A40	6720
x"00",	-- Hex Addr	1A41	6721
x"00",	-- Hex Addr	1A42	6722
x"00",	-- Hex Addr	1A43	6723
x"00",	-- Hex Addr	1A44	6724
x"00",	-- Hex Addr	1A45	6725
x"00",	-- Hex Addr	1A46	6726
x"00",	-- Hex Addr	1A47	6727
x"00",	-- Hex Addr	1A48	6728
x"00",	-- Hex Addr	1A49	6729
x"00",	-- Hex Addr	1A4A	6730
x"00",	-- Hex Addr	1A4B	6731
x"00",	-- Hex Addr	1A4C	6732
x"00",	-- Hex Addr	1A4D	6733
x"00",	-- Hex Addr	1A4E	6734
x"00",	-- Hex Addr	1A4F	6735
x"00",	-- Hex Addr	1A50	6736
x"00",	-- Hex Addr	1A51	6737
x"00",	-- Hex Addr	1A52	6738
x"00",	-- Hex Addr	1A53	6739
x"00",	-- Hex Addr	1A54	6740
x"00",	-- Hex Addr	1A55	6741
x"00",	-- Hex Addr	1A56	6742
x"00",	-- Hex Addr	1A57	6743
x"00",	-- Hex Addr	1A58	6744
x"00",	-- Hex Addr	1A59	6745
x"00",	-- Hex Addr	1A5A	6746
x"00",	-- Hex Addr	1A5B	6747
x"00",	-- Hex Addr	1A5C	6748
x"00",	-- Hex Addr	1A5D	6749
x"00",	-- Hex Addr	1A5E	6750
x"00",	-- Hex Addr	1A5F	6751
x"00",	-- Hex Addr	1A60	6752
x"00",	-- Hex Addr	1A61	6753
x"00",	-- Hex Addr	1A62	6754
x"00",	-- Hex Addr	1A63	6755
x"00",	-- Hex Addr	1A64	6756
x"00",	-- Hex Addr	1A65	6757
x"00",	-- Hex Addr	1A66	6758
x"00",	-- Hex Addr	1A67	6759
x"00",	-- Hex Addr	1A68	6760
x"00",	-- Hex Addr	1A69	6761
x"00",	-- Hex Addr	1A6A	6762
x"00",	-- Hex Addr	1A6B	6763
x"00",	-- Hex Addr	1A6C	6764
x"00",	-- Hex Addr	1A6D	6765
x"00",	-- Hex Addr	1A6E	6766
x"00",	-- Hex Addr	1A6F	6767
x"00",	-- Hex Addr	1A70	6768
x"00",	-- Hex Addr	1A71	6769
x"00",	-- Hex Addr	1A72	6770
x"00",	-- Hex Addr	1A73	6771
x"00",	-- Hex Addr	1A74	6772
x"00",	-- Hex Addr	1A75	6773
x"00",	-- Hex Addr	1A76	6774
x"00",	-- Hex Addr	1A77	6775
x"00",	-- Hex Addr	1A78	6776
x"00",	-- Hex Addr	1A79	6777
x"00",	-- Hex Addr	1A7A	6778
x"00",	-- Hex Addr	1A7B	6779
x"00",	-- Hex Addr	1A7C	6780
x"00",	-- Hex Addr	1A7D	6781
x"00",	-- Hex Addr	1A7E	6782
x"00",	-- Hex Addr	1A7F	6783
x"00",	-- Hex Addr	1A80	6784
x"00",	-- Hex Addr	1A81	6785
x"00",	-- Hex Addr	1A82	6786
x"00",	-- Hex Addr	1A83	6787
x"00",	-- Hex Addr	1A84	6788
x"00",	-- Hex Addr	1A85	6789
x"00",	-- Hex Addr	1A86	6790
x"00",	-- Hex Addr	1A87	6791
x"00",	-- Hex Addr	1A88	6792
x"00",	-- Hex Addr	1A89	6793
x"00",	-- Hex Addr	1A8A	6794
x"00",	-- Hex Addr	1A8B	6795
x"00",	-- Hex Addr	1A8C	6796
x"00",	-- Hex Addr	1A8D	6797
x"00",	-- Hex Addr	1A8E	6798
x"00",	-- Hex Addr	1A8F	6799
x"00",	-- Hex Addr	1A90	6800
x"00",	-- Hex Addr	1A91	6801
x"00",	-- Hex Addr	1A92	6802
x"00",	-- Hex Addr	1A93	6803
x"00",	-- Hex Addr	1A94	6804
x"00",	-- Hex Addr	1A95	6805
x"00",	-- Hex Addr	1A96	6806
x"00",	-- Hex Addr	1A97	6807
x"00",	-- Hex Addr	1A98	6808
x"00",	-- Hex Addr	1A99	6809
x"00",	-- Hex Addr	1A9A	6810
x"00",	-- Hex Addr	1A9B	6811
x"00",	-- Hex Addr	1A9C	6812
x"00",	-- Hex Addr	1A9D	6813
x"00",	-- Hex Addr	1A9E	6814
x"00",	-- Hex Addr	1A9F	6815
x"00",	-- Hex Addr	1AA0	6816
x"00",	-- Hex Addr	1AA1	6817
x"00",	-- Hex Addr	1AA2	6818
x"00",	-- Hex Addr	1AA3	6819
x"00",	-- Hex Addr	1AA4	6820
x"00",	-- Hex Addr	1AA5	6821
x"00",	-- Hex Addr	1AA6	6822
x"00",	-- Hex Addr	1AA7	6823
x"00",	-- Hex Addr	1AA8	6824
x"00",	-- Hex Addr	1AA9	6825
x"00",	-- Hex Addr	1AAA	6826
x"00",	-- Hex Addr	1AAB	6827
x"00",	-- Hex Addr	1AAC	6828
x"00",	-- Hex Addr	1AAD	6829
x"00",	-- Hex Addr	1AAE	6830
x"00",	-- Hex Addr	1AAF	6831
x"00",	-- Hex Addr	1AB0	6832
x"00",	-- Hex Addr	1AB1	6833
x"00",	-- Hex Addr	1AB2	6834
x"00",	-- Hex Addr	1AB3	6835
x"00",	-- Hex Addr	1AB4	6836
x"00",	-- Hex Addr	1AB5	6837
x"00",	-- Hex Addr	1AB6	6838
x"00",	-- Hex Addr	1AB7	6839
x"00",	-- Hex Addr	1AB8	6840
x"00",	-- Hex Addr	1AB9	6841
x"00",	-- Hex Addr	1ABA	6842
x"00",	-- Hex Addr	1ABB	6843
x"00",	-- Hex Addr	1ABC	6844
x"00",	-- Hex Addr	1ABD	6845
x"00",	-- Hex Addr	1ABE	6846
x"00",	-- Hex Addr	1ABF	6847
x"00",	-- Hex Addr	1AC0	6848
x"00",	-- Hex Addr	1AC1	6849
x"00",	-- Hex Addr	1AC2	6850
x"00",	-- Hex Addr	1AC3	6851
x"00",	-- Hex Addr	1AC4	6852
x"00",	-- Hex Addr	1AC5	6853
x"00",	-- Hex Addr	1AC6	6854
x"00",	-- Hex Addr	1AC7	6855
x"00",	-- Hex Addr	1AC8	6856
x"00",	-- Hex Addr	1AC9	6857
x"00",	-- Hex Addr	1ACA	6858
x"00",	-- Hex Addr	1ACB	6859
x"00",	-- Hex Addr	1ACC	6860
x"00",	-- Hex Addr	1ACD	6861
x"00",	-- Hex Addr	1ACE	6862
x"00",	-- Hex Addr	1ACF	6863
x"00",	-- Hex Addr	1AD0	6864
x"00",	-- Hex Addr	1AD1	6865
x"00",	-- Hex Addr	1AD2	6866
x"00",	-- Hex Addr	1AD3	6867
x"00",	-- Hex Addr	1AD4	6868
x"00",	-- Hex Addr	1AD5	6869
x"00",	-- Hex Addr	1AD6	6870
x"00",	-- Hex Addr	1AD7	6871
x"00",	-- Hex Addr	1AD8	6872
x"00",	-- Hex Addr	1AD9	6873
x"00",	-- Hex Addr	1ADA	6874
x"00",	-- Hex Addr	1ADB	6875
x"00",	-- Hex Addr	1ADC	6876
x"00",	-- Hex Addr	1ADD	6877
x"00",	-- Hex Addr	1ADE	6878
x"00",	-- Hex Addr	1ADF	6879
x"00",	-- Hex Addr	1AE0	6880
x"00",	-- Hex Addr	1AE1	6881
x"00",	-- Hex Addr	1AE2	6882
x"00",	-- Hex Addr	1AE3	6883
x"00",	-- Hex Addr	1AE4	6884
x"00",	-- Hex Addr	1AE5	6885
x"00",	-- Hex Addr	1AE6	6886
x"00",	-- Hex Addr	1AE7	6887
x"00",	-- Hex Addr	1AE8	6888
x"00",	-- Hex Addr	1AE9	6889
x"00",	-- Hex Addr	1AEA	6890
x"00",	-- Hex Addr	1AEB	6891
x"00",	-- Hex Addr	1AEC	6892
x"00",	-- Hex Addr	1AED	6893
x"00",	-- Hex Addr	1AEE	6894
x"00",	-- Hex Addr	1AEF	6895
x"00",	-- Hex Addr	1AF0	6896
x"00",	-- Hex Addr	1AF1	6897
x"00",	-- Hex Addr	1AF2	6898
x"00",	-- Hex Addr	1AF3	6899
x"00",	-- Hex Addr	1AF4	6900
x"00",	-- Hex Addr	1AF5	6901
x"00",	-- Hex Addr	1AF6	6902
x"00",	-- Hex Addr	1AF7	6903
x"00",	-- Hex Addr	1AF8	6904
x"00",	-- Hex Addr	1AF9	6905
x"00",	-- Hex Addr	1AFA	6906
x"00",	-- Hex Addr	1AFB	6907
x"00",	-- Hex Addr	1AFC	6908
x"00",	-- Hex Addr	1AFD	6909
x"00",	-- Hex Addr	1AFE	6910
x"00",	-- Hex Addr	1AFF	6911
x"00",	-- Hex Addr	1B00	6912
x"00",	-- Hex Addr	1B01	6913
x"00",	-- Hex Addr	1B02	6914
x"00",	-- Hex Addr	1B03	6915
x"00",	-- Hex Addr	1B04	6916
x"00",	-- Hex Addr	1B05	6917
x"00",	-- Hex Addr	1B06	6918
x"00",	-- Hex Addr	1B07	6919
x"00",	-- Hex Addr	1B08	6920
x"00",	-- Hex Addr	1B09	6921
x"00",	-- Hex Addr	1B0A	6922
x"00",	-- Hex Addr	1B0B	6923
x"00",	-- Hex Addr	1B0C	6924
x"00",	-- Hex Addr	1B0D	6925
x"00",	-- Hex Addr	1B0E	6926
x"00",	-- Hex Addr	1B0F	6927
x"00",	-- Hex Addr	1B10	6928
x"00",	-- Hex Addr	1B11	6929
x"00",	-- Hex Addr	1B12	6930
x"00",	-- Hex Addr	1B13	6931
x"00",	-- Hex Addr	1B14	6932
x"00",	-- Hex Addr	1B15	6933
x"00",	-- Hex Addr	1B16	6934
x"00",	-- Hex Addr	1B17	6935
x"00",	-- Hex Addr	1B18	6936
x"00",	-- Hex Addr	1B19	6937
x"00",	-- Hex Addr	1B1A	6938
x"00",	-- Hex Addr	1B1B	6939
x"00",	-- Hex Addr	1B1C	6940
x"00",	-- Hex Addr	1B1D	6941
x"00",	-- Hex Addr	1B1E	6942
x"00",	-- Hex Addr	1B1F	6943
x"00",	-- Hex Addr	1B20	6944
x"00",	-- Hex Addr	1B21	6945
x"00",	-- Hex Addr	1B22	6946
x"00",	-- Hex Addr	1B23	6947
x"00",	-- Hex Addr	1B24	6948
x"00",	-- Hex Addr	1B25	6949
x"00",	-- Hex Addr	1B26	6950
x"00",	-- Hex Addr	1B27	6951
x"00",	-- Hex Addr	1B28	6952
x"00",	-- Hex Addr	1B29	6953
x"00",	-- Hex Addr	1B2A	6954
x"00",	-- Hex Addr	1B2B	6955
x"00",	-- Hex Addr	1B2C	6956
x"00",	-- Hex Addr	1B2D	6957
x"00",	-- Hex Addr	1B2E	6958
x"00",	-- Hex Addr	1B2F	6959
x"00",	-- Hex Addr	1B30	6960
x"00",	-- Hex Addr	1B31	6961
x"00",	-- Hex Addr	1B32	6962
x"00",	-- Hex Addr	1B33	6963
x"00",	-- Hex Addr	1B34	6964
x"00",	-- Hex Addr	1B35	6965
x"00",	-- Hex Addr	1B36	6966
x"00",	-- Hex Addr	1B37	6967
x"00",	-- Hex Addr	1B38	6968
x"00",	-- Hex Addr	1B39	6969
x"00",	-- Hex Addr	1B3A	6970
x"00",	-- Hex Addr	1B3B	6971
x"00",	-- Hex Addr	1B3C	6972
x"00",	-- Hex Addr	1B3D	6973
x"00",	-- Hex Addr	1B3E	6974
x"00",	-- Hex Addr	1B3F	6975
x"00",	-- Hex Addr	1B40	6976
x"00",	-- Hex Addr	1B41	6977
x"00",	-- Hex Addr	1B42	6978
x"00",	-- Hex Addr	1B43	6979
x"00",	-- Hex Addr	1B44	6980
x"00",	-- Hex Addr	1B45	6981
x"00",	-- Hex Addr	1B46	6982
x"00",	-- Hex Addr	1B47	6983
x"00",	-- Hex Addr	1B48	6984
x"00",	-- Hex Addr	1B49	6985
x"00",	-- Hex Addr	1B4A	6986
x"00",	-- Hex Addr	1B4B	6987
x"00",	-- Hex Addr	1B4C	6988
x"00",	-- Hex Addr	1B4D	6989
x"00",	-- Hex Addr	1B4E	6990
x"00",	-- Hex Addr	1B4F	6991
x"00",	-- Hex Addr	1B50	6992
x"00",	-- Hex Addr	1B51	6993
x"00",	-- Hex Addr	1B52	6994
x"00",	-- Hex Addr	1B53	6995
x"00",	-- Hex Addr	1B54	6996
x"00",	-- Hex Addr	1B55	6997
x"00",	-- Hex Addr	1B56	6998
x"00",	-- Hex Addr	1B57	6999
x"00",	-- Hex Addr	1B58	7000
x"00",	-- Hex Addr	1B59	7001
x"00",	-- Hex Addr	1B5A	7002
x"00",	-- Hex Addr	1B5B	7003
x"00",	-- Hex Addr	1B5C	7004
x"00",	-- Hex Addr	1B5D	7005
x"00",	-- Hex Addr	1B5E	7006
x"00",	-- Hex Addr	1B5F	7007
x"00",	-- Hex Addr	1B60	7008
x"00",	-- Hex Addr	1B61	7009
x"00",	-- Hex Addr	1B62	7010
x"00",	-- Hex Addr	1B63	7011
x"00",	-- Hex Addr	1B64	7012
x"00",	-- Hex Addr	1B65	7013
x"00",	-- Hex Addr	1B66	7014
x"00",	-- Hex Addr	1B67	7015
x"00",	-- Hex Addr	1B68	7016
x"00",	-- Hex Addr	1B69	7017
x"00",	-- Hex Addr	1B6A	7018
x"00",	-- Hex Addr	1B6B	7019
x"00",	-- Hex Addr	1B6C	7020
x"00",	-- Hex Addr	1B6D	7021
x"00",	-- Hex Addr	1B6E	7022
x"00",	-- Hex Addr	1B6F	7023
x"00",	-- Hex Addr	1B70	7024
x"00",	-- Hex Addr	1B71	7025
x"00",	-- Hex Addr	1B72	7026
x"00",	-- Hex Addr	1B73	7027
x"00",	-- Hex Addr	1B74	7028
x"00",	-- Hex Addr	1B75	7029
x"00",	-- Hex Addr	1B76	7030
x"00",	-- Hex Addr	1B77	7031
x"00",	-- Hex Addr	1B78	7032
x"00",	-- Hex Addr	1B79	7033
x"00",	-- Hex Addr	1B7A	7034
x"00",	-- Hex Addr	1B7B	7035
x"00",	-- Hex Addr	1B7C	7036
x"00",	-- Hex Addr	1B7D	7037
x"00",	-- Hex Addr	1B7E	7038
x"00",	-- Hex Addr	1B7F	7039
x"00",	-- Hex Addr	1B80	7040
x"00",	-- Hex Addr	1B81	7041
x"00",	-- Hex Addr	1B82	7042
x"00",	-- Hex Addr	1B83	7043
x"00",	-- Hex Addr	1B84	7044
x"00",	-- Hex Addr	1B85	7045
x"00",	-- Hex Addr	1B86	7046
x"00",	-- Hex Addr	1B87	7047
x"00",	-- Hex Addr	1B88	7048
x"00",	-- Hex Addr	1B89	7049
x"00",	-- Hex Addr	1B8A	7050
x"00",	-- Hex Addr	1B8B	7051
x"00",	-- Hex Addr	1B8C	7052
x"00",	-- Hex Addr	1B8D	7053
x"00",	-- Hex Addr	1B8E	7054
x"00",	-- Hex Addr	1B8F	7055
x"00",	-- Hex Addr	1B90	7056
x"00",	-- Hex Addr	1B91	7057
x"00",	-- Hex Addr	1B92	7058
x"00",	-- Hex Addr	1B93	7059
x"00",	-- Hex Addr	1B94	7060
x"00",	-- Hex Addr	1B95	7061
x"00",	-- Hex Addr	1B96	7062
x"00",	-- Hex Addr	1B97	7063
x"00",	-- Hex Addr	1B98	7064
x"00",	-- Hex Addr	1B99	7065
x"00",	-- Hex Addr	1B9A	7066
x"00",	-- Hex Addr	1B9B	7067
x"00",	-- Hex Addr	1B9C	7068
x"00",	-- Hex Addr	1B9D	7069
x"00",	-- Hex Addr	1B9E	7070
x"00",	-- Hex Addr	1B9F	7071
x"00",	-- Hex Addr	1BA0	7072
x"00",	-- Hex Addr	1BA1	7073
x"00",	-- Hex Addr	1BA2	7074
x"00",	-- Hex Addr	1BA3	7075
x"00",	-- Hex Addr	1BA4	7076
x"00",	-- Hex Addr	1BA5	7077
x"00",	-- Hex Addr	1BA6	7078
x"00",	-- Hex Addr	1BA7	7079
x"00",	-- Hex Addr	1BA8	7080
x"00",	-- Hex Addr	1BA9	7081
x"00",	-- Hex Addr	1BAA	7082
x"00",	-- Hex Addr	1BAB	7083
x"00",	-- Hex Addr	1BAC	7084
x"00",	-- Hex Addr	1BAD	7085
x"00",	-- Hex Addr	1BAE	7086
x"00",	-- Hex Addr	1BAF	7087
x"00",	-- Hex Addr	1BB0	7088
x"00",	-- Hex Addr	1BB1	7089
x"00",	-- Hex Addr	1BB2	7090
x"00",	-- Hex Addr	1BB3	7091
x"00",	-- Hex Addr	1BB4	7092
x"00",	-- Hex Addr	1BB5	7093
x"00",	-- Hex Addr	1BB6	7094
x"00",	-- Hex Addr	1BB7	7095
x"00",	-- Hex Addr	1BB8	7096
x"00",	-- Hex Addr	1BB9	7097
x"00",	-- Hex Addr	1BBA	7098
x"00",	-- Hex Addr	1BBB	7099
x"00",	-- Hex Addr	1BBC	7100
x"00",	-- Hex Addr	1BBD	7101
x"00",	-- Hex Addr	1BBE	7102
x"00",	-- Hex Addr	1BBF	7103
x"00",	-- Hex Addr	1BC0	7104
x"00",	-- Hex Addr	1BC1	7105
x"00",	-- Hex Addr	1BC2	7106
x"00",	-- Hex Addr	1BC3	7107
x"00",	-- Hex Addr	1BC4	7108
x"00",	-- Hex Addr	1BC5	7109
x"00",	-- Hex Addr	1BC6	7110
x"00",	-- Hex Addr	1BC7	7111
x"00",	-- Hex Addr	1BC8	7112
x"00",	-- Hex Addr	1BC9	7113
x"00",	-- Hex Addr	1BCA	7114
x"00",	-- Hex Addr	1BCB	7115
x"00",	-- Hex Addr	1BCC	7116
x"00",	-- Hex Addr	1BCD	7117
x"00",	-- Hex Addr	1BCE	7118
x"00",	-- Hex Addr	1BCF	7119
x"00",	-- Hex Addr	1BD0	7120
x"00",	-- Hex Addr	1BD1	7121
x"00",	-- Hex Addr	1BD2	7122
x"00",	-- Hex Addr	1BD3	7123
x"00",	-- Hex Addr	1BD4	7124
x"00",	-- Hex Addr	1BD5	7125
x"00",	-- Hex Addr	1BD6	7126
x"00",	-- Hex Addr	1BD7	7127
x"00",	-- Hex Addr	1BD8	7128
x"00",	-- Hex Addr	1BD9	7129
x"00",	-- Hex Addr	1BDA	7130
x"00",	-- Hex Addr	1BDB	7131
x"00",	-- Hex Addr	1BDC	7132
x"00",	-- Hex Addr	1BDD	7133
x"00",	-- Hex Addr	1BDE	7134
x"00",	-- Hex Addr	1BDF	7135
x"00",	-- Hex Addr	1BE0	7136
x"00",	-- Hex Addr	1BE1	7137
x"00",	-- Hex Addr	1BE2	7138
x"00",	-- Hex Addr	1BE3	7139
x"00",	-- Hex Addr	1BE4	7140
x"00",	-- Hex Addr	1BE5	7141
x"00",	-- Hex Addr	1BE6	7142
x"00",	-- Hex Addr	1BE7	7143
x"00",	-- Hex Addr	1BE8	7144
x"00",	-- Hex Addr	1BE9	7145
x"00",	-- Hex Addr	1BEA	7146
x"00",	-- Hex Addr	1BEB	7147
x"00",	-- Hex Addr	1BEC	7148
x"00",	-- Hex Addr	1BED	7149
x"00",	-- Hex Addr	1BEE	7150
x"00",	-- Hex Addr	1BEF	7151
x"00",	-- Hex Addr	1BF0	7152
x"00",	-- Hex Addr	1BF1	7153
x"00",	-- Hex Addr	1BF2	7154
x"00",	-- Hex Addr	1BF3	7155
x"00",	-- Hex Addr	1BF4	7156
x"00",	-- Hex Addr	1BF5	7157
x"00",	-- Hex Addr	1BF6	7158
x"00",	-- Hex Addr	1BF7	7159
x"00",	-- Hex Addr	1BF8	7160
x"00",	-- Hex Addr	1BF9	7161
x"00",	-- Hex Addr	1BFA	7162
x"00",	-- Hex Addr	1BFB	7163
x"00",	-- Hex Addr	1BFC	7164
x"00",	-- Hex Addr	1BFD	7165
x"00",	-- Hex Addr	1BFE	7166
x"00",	-- Hex Addr	1BFF	7167
x"00",	-- Hex Addr	1C00	7168
x"00",	-- Hex Addr	1C01	7169
x"00",	-- Hex Addr	1C02	7170
x"00",	-- Hex Addr	1C03	7171
x"00",	-- Hex Addr	1C04	7172
x"00",	-- Hex Addr	1C05	7173
x"00",	-- Hex Addr	1C06	7174
x"00",	-- Hex Addr	1C07	7175
x"00",	-- Hex Addr	1C08	7176
x"00",	-- Hex Addr	1C09	7177
x"00",	-- Hex Addr	1C0A	7178
x"00",	-- Hex Addr	1C0B	7179
x"00",	-- Hex Addr	1C0C	7180
x"00",	-- Hex Addr	1C0D	7181
x"00",	-- Hex Addr	1C0E	7182
x"00",	-- Hex Addr	1C0F	7183
x"00",	-- Hex Addr	1C10	7184
x"00",	-- Hex Addr	1C11	7185
x"00",	-- Hex Addr	1C12	7186
x"00",	-- Hex Addr	1C13	7187
x"00",	-- Hex Addr	1C14	7188
x"00",	-- Hex Addr	1C15	7189
x"00",	-- Hex Addr	1C16	7190
x"00",	-- Hex Addr	1C17	7191
x"00",	-- Hex Addr	1C18	7192
x"00",	-- Hex Addr	1C19	7193
x"00",	-- Hex Addr	1C1A	7194
x"00",	-- Hex Addr	1C1B	7195
x"00",	-- Hex Addr	1C1C	7196
x"00",	-- Hex Addr	1C1D	7197
x"00",	-- Hex Addr	1C1E	7198
x"00",	-- Hex Addr	1C1F	7199
x"00",	-- Hex Addr	1C20	7200
x"00",	-- Hex Addr	1C21	7201
x"00",	-- Hex Addr	1C22	7202
x"00",	-- Hex Addr	1C23	7203
x"00",	-- Hex Addr	1C24	7204
x"00",	-- Hex Addr	1C25	7205
x"00",	-- Hex Addr	1C26	7206
x"00",	-- Hex Addr	1C27	7207
x"00",	-- Hex Addr	1C28	7208
x"00",	-- Hex Addr	1C29	7209
x"00",	-- Hex Addr	1C2A	7210
x"00",	-- Hex Addr	1C2B	7211
x"00",	-- Hex Addr	1C2C	7212
x"00",	-- Hex Addr	1C2D	7213
x"00",	-- Hex Addr	1C2E	7214
x"00",	-- Hex Addr	1C2F	7215
x"00",	-- Hex Addr	1C30	7216
x"00",	-- Hex Addr	1C31	7217
x"00",	-- Hex Addr	1C32	7218
x"00",	-- Hex Addr	1C33	7219
x"00",	-- Hex Addr	1C34	7220
x"00",	-- Hex Addr	1C35	7221
x"00",	-- Hex Addr	1C36	7222
x"00",	-- Hex Addr	1C37	7223
x"00",	-- Hex Addr	1C38	7224
x"00",	-- Hex Addr	1C39	7225
x"00",	-- Hex Addr	1C3A	7226
x"00",	-- Hex Addr	1C3B	7227
x"00",	-- Hex Addr	1C3C	7228
x"00",	-- Hex Addr	1C3D	7229
x"00",	-- Hex Addr	1C3E	7230
x"00",	-- Hex Addr	1C3F	7231
x"00",	-- Hex Addr	1C40	7232
x"00",	-- Hex Addr	1C41	7233
x"00",	-- Hex Addr	1C42	7234
x"00",	-- Hex Addr	1C43	7235
x"00",	-- Hex Addr	1C44	7236
x"00",	-- Hex Addr	1C45	7237
x"00",	-- Hex Addr	1C46	7238
x"00",	-- Hex Addr	1C47	7239
x"00",	-- Hex Addr	1C48	7240
x"00",	-- Hex Addr	1C49	7241
x"00",	-- Hex Addr	1C4A	7242
x"00",	-- Hex Addr	1C4B	7243
x"00",	-- Hex Addr	1C4C	7244
x"00",	-- Hex Addr	1C4D	7245
x"00",	-- Hex Addr	1C4E	7246
x"00",	-- Hex Addr	1C4F	7247
x"00",	-- Hex Addr	1C50	7248
x"00",	-- Hex Addr	1C51	7249
x"00",	-- Hex Addr	1C52	7250
x"00",	-- Hex Addr	1C53	7251
x"00",	-- Hex Addr	1C54	7252
x"00",	-- Hex Addr	1C55	7253
x"00",	-- Hex Addr	1C56	7254
x"00",	-- Hex Addr	1C57	7255
x"00",	-- Hex Addr	1C58	7256
x"00",	-- Hex Addr	1C59	7257
x"00",	-- Hex Addr	1C5A	7258
x"00",	-- Hex Addr	1C5B	7259
x"00",	-- Hex Addr	1C5C	7260
x"00",	-- Hex Addr	1C5D	7261
x"00",	-- Hex Addr	1C5E	7262
x"00",	-- Hex Addr	1C5F	7263
x"00",	-- Hex Addr	1C60	7264
x"00",	-- Hex Addr	1C61	7265
x"00",	-- Hex Addr	1C62	7266
x"00",	-- Hex Addr	1C63	7267
x"00",	-- Hex Addr	1C64	7268
x"00",	-- Hex Addr	1C65	7269
x"00",	-- Hex Addr	1C66	7270
x"00",	-- Hex Addr	1C67	7271
x"00",	-- Hex Addr	1C68	7272
x"00",	-- Hex Addr	1C69	7273
x"00",	-- Hex Addr	1C6A	7274
x"00",	-- Hex Addr	1C6B	7275
x"00",	-- Hex Addr	1C6C	7276
x"00",	-- Hex Addr	1C6D	7277
x"00",	-- Hex Addr	1C6E	7278
x"00",	-- Hex Addr	1C6F	7279
x"00",	-- Hex Addr	1C70	7280
x"00",	-- Hex Addr	1C71	7281
x"00",	-- Hex Addr	1C72	7282
x"00",	-- Hex Addr	1C73	7283
x"00",	-- Hex Addr	1C74	7284
x"00",	-- Hex Addr	1C75	7285
x"00",	-- Hex Addr	1C76	7286
x"00",	-- Hex Addr	1C77	7287
x"00",	-- Hex Addr	1C78	7288
x"00",	-- Hex Addr	1C79	7289
x"00",	-- Hex Addr	1C7A	7290
x"00",	-- Hex Addr	1C7B	7291
x"00",	-- Hex Addr	1C7C	7292
x"00",	-- Hex Addr	1C7D	7293
x"00",	-- Hex Addr	1C7E	7294
x"00",	-- Hex Addr	1C7F	7295
x"00",	-- Hex Addr	1C80	7296
x"00",	-- Hex Addr	1C81	7297
x"00",	-- Hex Addr	1C82	7298
x"00",	-- Hex Addr	1C83	7299
x"00",	-- Hex Addr	1C84	7300
x"00",	-- Hex Addr	1C85	7301
x"00",	-- Hex Addr	1C86	7302
x"00",	-- Hex Addr	1C87	7303
x"00",	-- Hex Addr	1C88	7304
x"00",	-- Hex Addr	1C89	7305
x"00",	-- Hex Addr	1C8A	7306
x"00",	-- Hex Addr	1C8B	7307
x"00",	-- Hex Addr	1C8C	7308
x"00",	-- Hex Addr	1C8D	7309
x"00",	-- Hex Addr	1C8E	7310
x"00",	-- Hex Addr	1C8F	7311
x"00",	-- Hex Addr	1C90	7312
x"00",	-- Hex Addr	1C91	7313
x"00",	-- Hex Addr	1C92	7314
x"00",	-- Hex Addr	1C93	7315
x"00",	-- Hex Addr	1C94	7316
x"00",	-- Hex Addr	1C95	7317
x"00",	-- Hex Addr	1C96	7318
x"00",	-- Hex Addr	1C97	7319
x"00",	-- Hex Addr	1C98	7320
x"00",	-- Hex Addr	1C99	7321
x"00",	-- Hex Addr	1C9A	7322
x"00",	-- Hex Addr	1C9B	7323
x"00",	-- Hex Addr	1C9C	7324
x"00",	-- Hex Addr	1C9D	7325
x"00",	-- Hex Addr	1C9E	7326
x"00",	-- Hex Addr	1C9F	7327
x"00",	-- Hex Addr	1CA0	7328
x"00",	-- Hex Addr	1CA1	7329
x"00",	-- Hex Addr	1CA2	7330
x"00",	-- Hex Addr	1CA3	7331
x"00",	-- Hex Addr	1CA4	7332
x"00",	-- Hex Addr	1CA5	7333
x"00",	-- Hex Addr	1CA6	7334
x"00",	-- Hex Addr	1CA7	7335
x"00",	-- Hex Addr	1CA8	7336
x"00",	-- Hex Addr	1CA9	7337
x"00",	-- Hex Addr	1CAA	7338
x"00",	-- Hex Addr	1CAB	7339
x"00",	-- Hex Addr	1CAC	7340
x"00",	-- Hex Addr	1CAD	7341
x"00",	-- Hex Addr	1CAE	7342
x"00",	-- Hex Addr	1CAF	7343
x"00",	-- Hex Addr	1CB0	7344
x"00",	-- Hex Addr	1CB1	7345
x"00",	-- Hex Addr	1CB2	7346
x"00",	-- Hex Addr	1CB3	7347
x"00",	-- Hex Addr	1CB4	7348
x"00",	-- Hex Addr	1CB5	7349
x"00",	-- Hex Addr	1CB6	7350
x"00",	-- Hex Addr	1CB7	7351
x"00",	-- Hex Addr	1CB8	7352
x"00",	-- Hex Addr	1CB9	7353
x"00",	-- Hex Addr	1CBA	7354
x"00",	-- Hex Addr	1CBB	7355
x"00",	-- Hex Addr	1CBC	7356
x"00",	-- Hex Addr	1CBD	7357
x"00",	-- Hex Addr	1CBE	7358
x"00",	-- Hex Addr	1CBF	7359
x"00",	-- Hex Addr	1CC0	7360
x"00",	-- Hex Addr	1CC1	7361
x"00",	-- Hex Addr	1CC2	7362
x"00",	-- Hex Addr	1CC3	7363
x"00",	-- Hex Addr	1CC4	7364
x"00",	-- Hex Addr	1CC5	7365
x"00",	-- Hex Addr	1CC6	7366
x"00",	-- Hex Addr	1CC7	7367
x"00",	-- Hex Addr	1CC8	7368
x"00",	-- Hex Addr	1CC9	7369
x"00",	-- Hex Addr	1CCA	7370
x"00",	-- Hex Addr	1CCB	7371
x"00",	-- Hex Addr	1CCC	7372
x"00",	-- Hex Addr	1CCD	7373
x"00",	-- Hex Addr	1CCE	7374
x"00",	-- Hex Addr	1CCF	7375
x"00",	-- Hex Addr	1CD0	7376
x"00",	-- Hex Addr	1CD1	7377
x"00",	-- Hex Addr	1CD2	7378
x"00",	-- Hex Addr	1CD3	7379
x"00",	-- Hex Addr	1CD4	7380
x"00",	-- Hex Addr	1CD5	7381
x"00",	-- Hex Addr	1CD6	7382
x"00",	-- Hex Addr	1CD7	7383
x"00",	-- Hex Addr	1CD8	7384
x"00",	-- Hex Addr	1CD9	7385
x"00",	-- Hex Addr	1CDA	7386
x"00",	-- Hex Addr	1CDB	7387
x"00",	-- Hex Addr	1CDC	7388
x"00",	-- Hex Addr	1CDD	7389
x"00",	-- Hex Addr	1CDE	7390
x"00",	-- Hex Addr	1CDF	7391
x"00",	-- Hex Addr	1CE0	7392
x"00",	-- Hex Addr	1CE1	7393
x"00",	-- Hex Addr	1CE2	7394
x"00",	-- Hex Addr	1CE3	7395
x"00",	-- Hex Addr	1CE4	7396
x"00",	-- Hex Addr	1CE5	7397
x"00",	-- Hex Addr	1CE6	7398
x"00",	-- Hex Addr	1CE7	7399
x"00",	-- Hex Addr	1CE8	7400
x"00",	-- Hex Addr	1CE9	7401
x"00",	-- Hex Addr	1CEA	7402
x"00",	-- Hex Addr	1CEB	7403
x"00",	-- Hex Addr	1CEC	7404
x"00",	-- Hex Addr	1CED	7405
x"00",	-- Hex Addr	1CEE	7406
x"00",	-- Hex Addr	1CEF	7407
x"00",	-- Hex Addr	1CF0	7408
x"00",	-- Hex Addr	1CF1	7409
x"00",	-- Hex Addr	1CF2	7410
x"00",	-- Hex Addr	1CF3	7411
x"00",	-- Hex Addr	1CF4	7412
x"00",	-- Hex Addr	1CF5	7413
x"00",	-- Hex Addr	1CF6	7414
x"00",	-- Hex Addr	1CF7	7415
x"00",	-- Hex Addr	1CF8	7416
x"00",	-- Hex Addr	1CF9	7417
x"00",	-- Hex Addr	1CFA	7418
x"00",	-- Hex Addr	1CFB	7419
x"00",	-- Hex Addr	1CFC	7420
x"00",	-- Hex Addr	1CFD	7421
x"00",	-- Hex Addr	1CFE	7422
x"00",	-- Hex Addr	1CFF	7423
x"00",	-- Hex Addr	1D00	7424
x"00",	-- Hex Addr	1D01	7425
x"00",	-- Hex Addr	1D02	7426
x"00",	-- Hex Addr	1D03	7427
x"00",	-- Hex Addr	1D04	7428
x"00",	-- Hex Addr	1D05	7429
x"00",	-- Hex Addr	1D06	7430
x"00",	-- Hex Addr	1D07	7431
x"00",	-- Hex Addr	1D08	7432
x"00",	-- Hex Addr	1D09	7433
x"00",	-- Hex Addr	1D0A	7434
x"00",	-- Hex Addr	1D0B	7435
x"00",	-- Hex Addr	1D0C	7436
x"00",	-- Hex Addr	1D0D	7437
x"00",	-- Hex Addr	1D0E	7438
x"00",	-- Hex Addr	1D0F	7439
x"00",	-- Hex Addr	1D10	7440
x"00",	-- Hex Addr	1D11	7441
x"00",	-- Hex Addr	1D12	7442
x"00",	-- Hex Addr	1D13	7443
x"00",	-- Hex Addr	1D14	7444
x"00",	-- Hex Addr	1D15	7445
x"00",	-- Hex Addr	1D16	7446
x"00",	-- Hex Addr	1D17	7447
x"00",	-- Hex Addr	1D18	7448
x"00",	-- Hex Addr	1D19	7449
x"00",	-- Hex Addr	1D1A	7450
x"00",	-- Hex Addr	1D1B	7451
x"00",	-- Hex Addr	1D1C	7452
x"00",	-- Hex Addr	1D1D	7453
x"00",	-- Hex Addr	1D1E	7454
x"00",	-- Hex Addr	1D1F	7455
x"00",	-- Hex Addr	1D20	7456
x"00",	-- Hex Addr	1D21	7457
x"00",	-- Hex Addr	1D22	7458
x"00",	-- Hex Addr	1D23	7459
x"00",	-- Hex Addr	1D24	7460
x"00",	-- Hex Addr	1D25	7461
x"00",	-- Hex Addr	1D26	7462
x"00",	-- Hex Addr	1D27	7463
x"00",	-- Hex Addr	1D28	7464
x"00",	-- Hex Addr	1D29	7465
x"00",	-- Hex Addr	1D2A	7466
x"00",	-- Hex Addr	1D2B	7467
x"00",	-- Hex Addr	1D2C	7468
x"00",	-- Hex Addr	1D2D	7469
x"00",	-- Hex Addr	1D2E	7470
x"00",	-- Hex Addr	1D2F	7471
x"00",	-- Hex Addr	1D30	7472
x"00",	-- Hex Addr	1D31	7473
x"00",	-- Hex Addr	1D32	7474
x"00",	-- Hex Addr	1D33	7475
x"00",	-- Hex Addr	1D34	7476
x"00",	-- Hex Addr	1D35	7477
x"00",	-- Hex Addr	1D36	7478
x"00",	-- Hex Addr	1D37	7479
x"00",	-- Hex Addr	1D38	7480
x"00",	-- Hex Addr	1D39	7481
x"00",	-- Hex Addr	1D3A	7482
x"00",	-- Hex Addr	1D3B	7483
x"00",	-- Hex Addr	1D3C	7484
x"00",	-- Hex Addr	1D3D	7485
x"00",	-- Hex Addr	1D3E	7486
x"00",	-- Hex Addr	1D3F	7487
x"00",	-- Hex Addr	1D40	7488
x"00",	-- Hex Addr	1D41	7489
x"00",	-- Hex Addr	1D42	7490
x"00",	-- Hex Addr	1D43	7491
x"00",	-- Hex Addr	1D44	7492
x"00",	-- Hex Addr	1D45	7493
x"00",	-- Hex Addr	1D46	7494
x"00",	-- Hex Addr	1D47	7495
x"00",	-- Hex Addr	1D48	7496
x"00",	-- Hex Addr	1D49	7497
x"00",	-- Hex Addr	1D4A	7498
x"00",	-- Hex Addr	1D4B	7499
x"00",	-- Hex Addr	1D4C	7500
x"00",	-- Hex Addr	1D4D	7501
x"00",	-- Hex Addr	1D4E	7502
x"00",	-- Hex Addr	1D4F	7503
x"00",	-- Hex Addr	1D50	7504
x"00",	-- Hex Addr	1D51	7505
x"00",	-- Hex Addr	1D52	7506
x"00",	-- Hex Addr	1D53	7507
x"00",	-- Hex Addr	1D54	7508
x"00",	-- Hex Addr	1D55	7509
x"00",	-- Hex Addr	1D56	7510
x"00",	-- Hex Addr	1D57	7511
x"00",	-- Hex Addr	1D58	7512
x"00",	-- Hex Addr	1D59	7513
x"00",	-- Hex Addr	1D5A	7514
x"00",	-- Hex Addr	1D5B	7515
x"00",	-- Hex Addr	1D5C	7516
x"00",	-- Hex Addr	1D5D	7517
x"00",	-- Hex Addr	1D5E	7518
x"00",	-- Hex Addr	1D5F	7519
x"00",	-- Hex Addr	1D60	7520
x"00",	-- Hex Addr	1D61	7521
x"00",	-- Hex Addr	1D62	7522
x"00",	-- Hex Addr	1D63	7523
x"00",	-- Hex Addr	1D64	7524
x"00",	-- Hex Addr	1D65	7525
x"00",	-- Hex Addr	1D66	7526
x"00",	-- Hex Addr	1D67	7527
x"00",	-- Hex Addr	1D68	7528
x"00",	-- Hex Addr	1D69	7529
x"00",	-- Hex Addr	1D6A	7530
x"00",	-- Hex Addr	1D6B	7531
x"00",	-- Hex Addr	1D6C	7532
x"00",	-- Hex Addr	1D6D	7533
x"00",	-- Hex Addr	1D6E	7534
x"00",	-- Hex Addr	1D6F	7535
x"00",	-- Hex Addr	1D70	7536
x"00",	-- Hex Addr	1D71	7537
x"00",	-- Hex Addr	1D72	7538
x"00",	-- Hex Addr	1D73	7539
x"00",	-- Hex Addr	1D74	7540
x"00",	-- Hex Addr	1D75	7541
x"00",	-- Hex Addr	1D76	7542
x"00",	-- Hex Addr	1D77	7543
x"00",	-- Hex Addr	1D78	7544
x"00",	-- Hex Addr	1D79	7545
x"00",	-- Hex Addr	1D7A	7546
x"00",	-- Hex Addr	1D7B	7547
x"00",	-- Hex Addr	1D7C	7548
x"00",	-- Hex Addr	1D7D	7549
x"00",	-- Hex Addr	1D7E	7550
x"00",	-- Hex Addr	1D7F	7551
x"00",	-- Hex Addr	1D80	7552
x"00",	-- Hex Addr	1D81	7553
x"00",	-- Hex Addr	1D82	7554
x"00",	-- Hex Addr	1D83	7555
x"00",	-- Hex Addr	1D84	7556
x"00",	-- Hex Addr	1D85	7557
x"00",	-- Hex Addr	1D86	7558
x"00",	-- Hex Addr	1D87	7559
x"00",	-- Hex Addr	1D88	7560
x"00",	-- Hex Addr	1D89	7561
x"00",	-- Hex Addr	1D8A	7562
x"00",	-- Hex Addr	1D8B	7563
x"00",	-- Hex Addr	1D8C	7564
x"00",	-- Hex Addr	1D8D	7565
x"00",	-- Hex Addr	1D8E	7566
x"00",	-- Hex Addr	1D8F	7567
x"00",	-- Hex Addr	1D90	7568
x"00",	-- Hex Addr	1D91	7569
x"00",	-- Hex Addr	1D92	7570
x"00",	-- Hex Addr	1D93	7571
x"00",	-- Hex Addr	1D94	7572
x"00",	-- Hex Addr	1D95	7573
x"00",	-- Hex Addr	1D96	7574
x"00",	-- Hex Addr	1D97	7575
x"00",	-- Hex Addr	1D98	7576
x"00",	-- Hex Addr	1D99	7577
x"00",	-- Hex Addr	1D9A	7578
x"00",	-- Hex Addr	1D9B	7579
x"00",	-- Hex Addr	1D9C	7580
x"00",	-- Hex Addr	1D9D	7581
x"00",	-- Hex Addr	1D9E	7582
x"00",	-- Hex Addr	1D9F	7583
x"00",	-- Hex Addr	1DA0	7584
x"00",	-- Hex Addr	1DA1	7585
x"00",	-- Hex Addr	1DA2	7586
x"00",	-- Hex Addr	1DA3	7587
x"00",	-- Hex Addr	1DA4	7588
x"00",	-- Hex Addr	1DA5	7589
x"00",	-- Hex Addr	1DA6	7590
x"00",	-- Hex Addr	1DA7	7591
x"00",	-- Hex Addr	1DA8	7592
x"00",	-- Hex Addr	1DA9	7593
x"00",	-- Hex Addr	1DAA	7594
x"00",	-- Hex Addr	1DAB	7595
x"00",	-- Hex Addr	1DAC	7596
x"00",	-- Hex Addr	1DAD	7597
x"00",	-- Hex Addr	1DAE	7598
x"00",	-- Hex Addr	1DAF	7599
x"00",	-- Hex Addr	1DB0	7600
x"00",	-- Hex Addr	1DB1	7601
x"00",	-- Hex Addr	1DB2	7602
x"00",	-- Hex Addr	1DB3	7603
x"00",	-- Hex Addr	1DB4	7604
x"00",	-- Hex Addr	1DB5	7605
x"00",	-- Hex Addr	1DB6	7606
x"00",	-- Hex Addr	1DB7	7607
x"00",	-- Hex Addr	1DB8	7608
x"00",	-- Hex Addr	1DB9	7609
x"00",	-- Hex Addr	1DBA	7610
x"00",	-- Hex Addr	1DBB	7611
x"00",	-- Hex Addr	1DBC	7612
x"00",	-- Hex Addr	1DBD	7613
x"00",	-- Hex Addr	1DBE	7614
x"00",	-- Hex Addr	1DBF	7615
x"00",	-- Hex Addr	1DC0	7616
x"00",	-- Hex Addr	1DC1	7617
x"00",	-- Hex Addr	1DC2	7618
x"00",	-- Hex Addr	1DC3	7619
x"00",	-- Hex Addr	1DC4	7620
x"00",	-- Hex Addr	1DC5	7621
x"00",	-- Hex Addr	1DC6	7622
x"00",	-- Hex Addr	1DC7	7623
x"00",	-- Hex Addr	1DC8	7624
x"00",	-- Hex Addr	1DC9	7625
x"00",	-- Hex Addr	1DCA	7626
x"00",	-- Hex Addr	1DCB	7627
x"00",	-- Hex Addr	1DCC	7628
x"00",	-- Hex Addr	1DCD	7629
x"00",	-- Hex Addr	1DCE	7630
x"00",	-- Hex Addr	1DCF	7631
x"00",	-- Hex Addr	1DD0	7632
x"00",	-- Hex Addr	1DD1	7633
x"00",	-- Hex Addr	1DD2	7634
x"00",	-- Hex Addr	1DD3	7635
x"00",	-- Hex Addr	1DD4	7636
x"00",	-- Hex Addr	1DD5	7637
x"00",	-- Hex Addr	1DD6	7638
x"00",	-- Hex Addr	1DD7	7639
x"00",	-- Hex Addr	1DD8	7640
x"00",	-- Hex Addr	1DD9	7641
x"00",	-- Hex Addr	1DDA	7642
x"00",	-- Hex Addr	1DDB	7643
x"00",	-- Hex Addr	1DDC	7644
x"00",	-- Hex Addr	1DDD	7645
x"00",	-- Hex Addr	1DDE	7646
x"00",	-- Hex Addr	1DDF	7647
x"00",	-- Hex Addr	1DE0	7648
x"00",	-- Hex Addr	1DE1	7649
x"00",	-- Hex Addr	1DE2	7650
x"00",	-- Hex Addr	1DE3	7651
x"00",	-- Hex Addr	1DE4	7652
x"00",	-- Hex Addr	1DE5	7653
x"00",	-- Hex Addr	1DE6	7654
x"00",	-- Hex Addr	1DE7	7655
x"00",	-- Hex Addr	1DE8	7656
x"00",	-- Hex Addr	1DE9	7657
x"00",	-- Hex Addr	1DEA	7658
x"00",	-- Hex Addr	1DEB	7659
x"00",	-- Hex Addr	1DEC	7660
x"00",	-- Hex Addr	1DED	7661
x"00",	-- Hex Addr	1DEE	7662
x"00",	-- Hex Addr	1DEF	7663
x"00",	-- Hex Addr	1DF0	7664
x"00",	-- Hex Addr	1DF1	7665
x"00",	-- Hex Addr	1DF2	7666
x"00",	-- Hex Addr	1DF3	7667
x"00",	-- Hex Addr	1DF4	7668
x"00",	-- Hex Addr	1DF5	7669
x"00",	-- Hex Addr	1DF6	7670
x"00",	-- Hex Addr	1DF7	7671
x"00",	-- Hex Addr	1DF8	7672
x"00",	-- Hex Addr	1DF9	7673
x"00",	-- Hex Addr	1DFA	7674
x"00",	-- Hex Addr	1DFB	7675
x"00",	-- Hex Addr	1DFC	7676
x"00",	-- Hex Addr	1DFD	7677
x"00",	-- Hex Addr	1DFE	7678
x"00",	-- Hex Addr	1DFF	7679
x"00",	-- Hex Addr	1E00	7680
x"00",	-- Hex Addr	1E01	7681
x"00",	-- Hex Addr	1E02	7682
x"00",	-- Hex Addr	1E03	7683
x"00",	-- Hex Addr	1E04	7684
x"00",	-- Hex Addr	1E05	7685
x"00",	-- Hex Addr	1E06	7686
x"00",	-- Hex Addr	1E07	7687
x"00",	-- Hex Addr	1E08	7688
x"00",	-- Hex Addr	1E09	7689
x"00",	-- Hex Addr	1E0A	7690
x"00",	-- Hex Addr	1E0B	7691
x"00",	-- Hex Addr	1E0C	7692
x"00",	-- Hex Addr	1E0D	7693
x"00",	-- Hex Addr	1E0E	7694
x"00",	-- Hex Addr	1E0F	7695
x"00",	-- Hex Addr	1E10	7696
x"00",	-- Hex Addr	1E11	7697
x"00",	-- Hex Addr	1E12	7698
x"00",	-- Hex Addr	1E13	7699
x"00",	-- Hex Addr	1E14	7700
x"00",	-- Hex Addr	1E15	7701
x"00",	-- Hex Addr	1E16	7702
x"00",	-- Hex Addr	1E17	7703
x"00",	-- Hex Addr	1E18	7704
x"00",	-- Hex Addr	1E19	7705
x"00",	-- Hex Addr	1E1A	7706
x"00",	-- Hex Addr	1E1B	7707
x"00",	-- Hex Addr	1E1C	7708
x"00",	-- Hex Addr	1E1D	7709
x"00",	-- Hex Addr	1E1E	7710
x"00",	-- Hex Addr	1E1F	7711
x"00",	-- Hex Addr	1E20	7712
x"00",	-- Hex Addr	1E21	7713
x"00",	-- Hex Addr	1E22	7714
x"00",	-- Hex Addr	1E23	7715
x"00",	-- Hex Addr	1E24	7716
x"00",	-- Hex Addr	1E25	7717
x"00",	-- Hex Addr	1E26	7718
x"00",	-- Hex Addr	1E27	7719
x"00",	-- Hex Addr	1E28	7720
x"00",	-- Hex Addr	1E29	7721
x"00",	-- Hex Addr	1E2A	7722
x"00",	-- Hex Addr	1E2B	7723
x"00",	-- Hex Addr	1E2C	7724
x"00",	-- Hex Addr	1E2D	7725
x"00",	-- Hex Addr	1E2E	7726
x"00",	-- Hex Addr	1E2F	7727
x"00",	-- Hex Addr	1E30	7728
x"00",	-- Hex Addr	1E31	7729
x"00",	-- Hex Addr	1E32	7730
x"00",	-- Hex Addr	1E33	7731
x"00",	-- Hex Addr	1E34	7732
x"00",	-- Hex Addr	1E35	7733
x"00",	-- Hex Addr	1E36	7734
x"00",	-- Hex Addr	1E37	7735
x"00",	-- Hex Addr	1E38	7736
x"00",	-- Hex Addr	1E39	7737
x"00",	-- Hex Addr	1E3A	7738
x"00",	-- Hex Addr	1E3B	7739
x"00",	-- Hex Addr	1E3C	7740
x"00",	-- Hex Addr	1E3D	7741
x"00",	-- Hex Addr	1E3E	7742
x"00",	-- Hex Addr	1E3F	7743
x"00",	-- Hex Addr	1E40	7744
x"00",	-- Hex Addr	1E41	7745
x"00",	-- Hex Addr	1E42	7746
x"00",	-- Hex Addr	1E43	7747
x"00",	-- Hex Addr	1E44	7748
x"00",	-- Hex Addr	1E45	7749
x"00",	-- Hex Addr	1E46	7750
x"00",	-- Hex Addr	1E47	7751
x"00",	-- Hex Addr	1E48	7752
x"00",	-- Hex Addr	1E49	7753
x"00",	-- Hex Addr	1E4A	7754
x"00",	-- Hex Addr	1E4B	7755
x"00",	-- Hex Addr	1E4C	7756
x"00",	-- Hex Addr	1E4D	7757
x"00",	-- Hex Addr	1E4E	7758
x"00",	-- Hex Addr	1E4F	7759
x"00",	-- Hex Addr	1E50	7760
x"00",	-- Hex Addr	1E51	7761
x"00",	-- Hex Addr	1E52	7762
x"00",	-- Hex Addr	1E53	7763
x"00",	-- Hex Addr	1E54	7764
x"00",	-- Hex Addr	1E55	7765
x"00",	-- Hex Addr	1E56	7766
x"00",	-- Hex Addr	1E57	7767
x"00",	-- Hex Addr	1E58	7768
x"00",	-- Hex Addr	1E59	7769
x"00",	-- Hex Addr	1E5A	7770
x"00",	-- Hex Addr	1E5B	7771
x"00",	-- Hex Addr	1E5C	7772
x"00",	-- Hex Addr	1E5D	7773
x"00",	-- Hex Addr	1E5E	7774
x"00",	-- Hex Addr	1E5F	7775
x"00",	-- Hex Addr	1E60	7776
x"00",	-- Hex Addr	1E61	7777
x"00",	-- Hex Addr	1E62	7778
x"00",	-- Hex Addr	1E63	7779
x"00",	-- Hex Addr	1E64	7780
x"00",	-- Hex Addr	1E65	7781
x"00",	-- Hex Addr	1E66	7782
x"00",	-- Hex Addr	1E67	7783
x"00",	-- Hex Addr	1E68	7784
x"00",	-- Hex Addr	1E69	7785
x"00",	-- Hex Addr	1E6A	7786
x"00",	-- Hex Addr	1E6B	7787
x"00",	-- Hex Addr	1E6C	7788
x"00",	-- Hex Addr	1E6D	7789
x"00",	-- Hex Addr	1E6E	7790
x"00",	-- Hex Addr	1E6F	7791
x"00",	-- Hex Addr	1E70	7792
x"00",	-- Hex Addr	1E71	7793
x"00",	-- Hex Addr	1E72	7794
x"00",	-- Hex Addr	1E73	7795
x"00",	-- Hex Addr	1E74	7796
x"00",	-- Hex Addr	1E75	7797
x"00",	-- Hex Addr	1E76	7798
x"00",	-- Hex Addr	1E77	7799
x"00",	-- Hex Addr	1E78	7800
x"00",	-- Hex Addr	1E79	7801
x"00",	-- Hex Addr	1E7A	7802
x"00",	-- Hex Addr	1E7B	7803
x"00",	-- Hex Addr	1E7C	7804
x"00",	-- Hex Addr	1E7D	7805
x"00",	-- Hex Addr	1E7E	7806
x"00",	-- Hex Addr	1E7F	7807
x"00",	-- Hex Addr	1E80	7808
x"00",	-- Hex Addr	1E81	7809
x"00",	-- Hex Addr	1E82	7810
x"00",	-- Hex Addr	1E83	7811
x"00",	-- Hex Addr	1E84	7812
x"00",	-- Hex Addr	1E85	7813
x"00",	-- Hex Addr	1E86	7814
x"00",	-- Hex Addr	1E87	7815
x"00",	-- Hex Addr	1E88	7816
x"00",	-- Hex Addr	1E89	7817
x"00",	-- Hex Addr	1E8A	7818
x"00",	-- Hex Addr	1E8B	7819
x"00",	-- Hex Addr	1E8C	7820
x"00",	-- Hex Addr	1E8D	7821
x"00",	-- Hex Addr	1E8E	7822
x"00",	-- Hex Addr	1E8F	7823
x"00",	-- Hex Addr	1E90	7824
x"00",	-- Hex Addr	1E91	7825
x"00",	-- Hex Addr	1E92	7826
x"00",	-- Hex Addr	1E93	7827
x"00",	-- Hex Addr	1E94	7828
x"00",	-- Hex Addr	1E95	7829
x"00",	-- Hex Addr	1E96	7830
x"00",	-- Hex Addr	1E97	7831
x"00",	-- Hex Addr	1E98	7832
x"00",	-- Hex Addr	1E99	7833
x"00",	-- Hex Addr	1E9A	7834
x"00",	-- Hex Addr	1E9B	7835
x"00",	-- Hex Addr	1E9C	7836
x"00",	-- Hex Addr	1E9D	7837
x"00",	-- Hex Addr	1E9E	7838
x"00",	-- Hex Addr	1E9F	7839
x"00",	-- Hex Addr	1EA0	7840
x"00",	-- Hex Addr	1EA1	7841
x"00",	-- Hex Addr	1EA2	7842
x"00",	-- Hex Addr	1EA3	7843
x"00",	-- Hex Addr	1EA4	7844
x"00",	-- Hex Addr	1EA5	7845
x"00",	-- Hex Addr	1EA6	7846
x"00",	-- Hex Addr	1EA7	7847
x"00",	-- Hex Addr	1EA8	7848
x"00",	-- Hex Addr	1EA9	7849
x"00",	-- Hex Addr	1EAA	7850
x"00",	-- Hex Addr	1EAB	7851
x"00",	-- Hex Addr	1EAC	7852
x"00",	-- Hex Addr	1EAD	7853
x"00",	-- Hex Addr	1EAE	7854
x"00",	-- Hex Addr	1EAF	7855
x"00",	-- Hex Addr	1EB0	7856
x"00",	-- Hex Addr	1EB1	7857
x"00",	-- Hex Addr	1EB2	7858
x"00",	-- Hex Addr	1EB3	7859
x"00",	-- Hex Addr	1EB4	7860
x"00",	-- Hex Addr	1EB5	7861
x"00",	-- Hex Addr	1EB6	7862
x"00",	-- Hex Addr	1EB7	7863
x"00",	-- Hex Addr	1EB8	7864
x"00",	-- Hex Addr	1EB9	7865
x"00",	-- Hex Addr	1EBA	7866
x"00",	-- Hex Addr	1EBB	7867
x"00",	-- Hex Addr	1EBC	7868
x"00",	-- Hex Addr	1EBD	7869
x"00",	-- Hex Addr	1EBE	7870
x"00",	-- Hex Addr	1EBF	7871
x"00",	-- Hex Addr	1EC0	7872
x"00",	-- Hex Addr	1EC1	7873
x"00",	-- Hex Addr	1EC2	7874
x"00",	-- Hex Addr	1EC3	7875
x"00",	-- Hex Addr	1EC4	7876
x"00",	-- Hex Addr	1EC5	7877
x"00",	-- Hex Addr	1EC6	7878
x"00",	-- Hex Addr	1EC7	7879
x"00",	-- Hex Addr	1EC8	7880
x"00",	-- Hex Addr	1EC9	7881
x"00",	-- Hex Addr	1ECA	7882
x"00",	-- Hex Addr	1ECB	7883
x"00",	-- Hex Addr	1ECC	7884
x"00",	-- Hex Addr	1ECD	7885
x"00",	-- Hex Addr	1ECE	7886
x"00",	-- Hex Addr	1ECF	7887
x"00",	-- Hex Addr	1ED0	7888
x"00",	-- Hex Addr	1ED1	7889
x"00",	-- Hex Addr	1ED2	7890
x"00",	-- Hex Addr	1ED3	7891
x"00",	-- Hex Addr	1ED4	7892
x"00",	-- Hex Addr	1ED5	7893
x"00",	-- Hex Addr	1ED6	7894
x"00",	-- Hex Addr	1ED7	7895
x"00",	-- Hex Addr	1ED8	7896
x"00",	-- Hex Addr	1ED9	7897
x"00",	-- Hex Addr	1EDA	7898
x"00",	-- Hex Addr	1EDB	7899
x"00",	-- Hex Addr	1EDC	7900
x"00",	-- Hex Addr	1EDD	7901
x"00",	-- Hex Addr	1EDE	7902
x"00",	-- Hex Addr	1EDF	7903
x"00",	-- Hex Addr	1EE0	7904
x"00",	-- Hex Addr	1EE1	7905
x"00",	-- Hex Addr	1EE2	7906
x"00",	-- Hex Addr	1EE3	7907
x"00",	-- Hex Addr	1EE4	7908
x"00",	-- Hex Addr	1EE5	7909
x"00",	-- Hex Addr	1EE6	7910
x"00",	-- Hex Addr	1EE7	7911
x"00",	-- Hex Addr	1EE8	7912
x"00",	-- Hex Addr	1EE9	7913
x"00",	-- Hex Addr	1EEA	7914
x"00",	-- Hex Addr	1EEB	7915
x"00",	-- Hex Addr	1EEC	7916
x"00",	-- Hex Addr	1EED	7917
x"00",	-- Hex Addr	1EEE	7918
x"00",	-- Hex Addr	1EEF	7919
x"00",	-- Hex Addr	1EF0	7920
x"00",	-- Hex Addr	1EF1	7921
x"00",	-- Hex Addr	1EF2	7922
x"00",	-- Hex Addr	1EF3	7923
x"00",	-- Hex Addr	1EF4	7924
x"00",	-- Hex Addr	1EF5	7925
x"00",	-- Hex Addr	1EF6	7926
x"00",	-- Hex Addr	1EF7	7927
x"00",	-- Hex Addr	1EF8	7928
x"00",	-- Hex Addr	1EF9	7929
x"00",	-- Hex Addr	1EFA	7930
x"00",	-- Hex Addr	1EFB	7931
x"00",	-- Hex Addr	1EFC	7932
x"00",	-- Hex Addr	1EFD	7933
x"00",	-- Hex Addr	1EFE	7934
x"00",	-- Hex Addr	1EFF	7935
x"00",	-- Hex Addr	1F00	7936
x"00",	-- Hex Addr	1F01	7937
x"00",	-- Hex Addr	1F02	7938
x"00",	-- Hex Addr	1F03	7939
x"00",	-- Hex Addr	1F04	7940
x"00",	-- Hex Addr	1F05	7941
x"00",	-- Hex Addr	1F06	7942
x"00",	-- Hex Addr	1F07	7943
x"00",	-- Hex Addr	1F08	7944
x"00",	-- Hex Addr	1F09	7945
x"00",	-- Hex Addr	1F0A	7946
x"00",	-- Hex Addr	1F0B	7947
x"00",	-- Hex Addr	1F0C	7948
x"00",	-- Hex Addr	1F0D	7949
x"00",	-- Hex Addr	1F0E	7950
x"00",	-- Hex Addr	1F0F	7951
x"00",	-- Hex Addr	1F10	7952
x"00",	-- Hex Addr	1F11	7953
x"00",	-- Hex Addr	1F12	7954
x"00",	-- Hex Addr	1F13	7955
x"00",	-- Hex Addr	1F14	7956
x"00",	-- Hex Addr	1F15	7957
x"00",	-- Hex Addr	1F16	7958
x"00",	-- Hex Addr	1F17	7959
x"00",	-- Hex Addr	1F18	7960
x"00",	-- Hex Addr	1F19	7961
x"00",	-- Hex Addr	1F1A	7962
x"00",	-- Hex Addr	1F1B	7963
x"00",	-- Hex Addr	1F1C	7964
x"00",	-- Hex Addr	1F1D	7965
x"00",	-- Hex Addr	1F1E	7966
x"00",	-- Hex Addr	1F1F	7967
x"00",	-- Hex Addr	1F20	7968
x"00",	-- Hex Addr	1F21	7969
x"00",	-- Hex Addr	1F22	7970
x"00",	-- Hex Addr	1F23	7971
x"00",	-- Hex Addr	1F24	7972
x"00",	-- Hex Addr	1F25	7973
x"00",	-- Hex Addr	1F26	7974
x"00",	-- Hex Addr	1F27	7975
x"00",	-- Hex Addr	1F28	7976
x"00",	-- Hex Addr	1F29	7977
x"00",	-- Hex Addr	1F2A	7978
x"00",	-- Hex Addr	1F2B	7979
x"00",	-- Hex Addr	1F2C	7980
x"00",	-- Hex Addr	1F2D	7981
x"00",	-- Hex Addr	1F2E	7982
x"00",	-- Hex Addr	1F2F	7983
x"00",	-- Hex Addr	1F30	7984
x"00",	-- Hex Addr	1F31	7985
x"00",	-- Hex Addr	1F32	7986
x"00",	-- Hex Addr	1F33	7987
x"00",	-- Hex Addr	1F34	7988
x"00",	-- Hex Addr	1F35	7989
x"00",	-- Hex Addr	1F36	7990
x"00",	-- Hex Addr	1F37	7991
x"00",	-- Hex Addr	1F38	7992
x"00",	-- Hex Addr	1F39	7993
x"00",	-- Hex Addr	1F3A	7994
x"00",	-- Hex Addr	1F3B	7995
x"00",	-- Hex Addr	1F3C	7996
x"00",	-- Hex Addr	1F3D	7997
x"00",	-- Hex Addr	1F3E	7998
x"00",	-- Hex Addr	1F3F	7999
x"00",	-- Hex Addr	1F40	8000
x"00",	-- Hex Addr	1F41	8001
x"00",	-- Hex Addr	1F42	8002
x"00",	-- Hex Addr	1F43	8003
x"00",	-- Hex Addr	1F44	8004
x"00",	-- Hex Addr	1F45	8005
x"00",	-- Hex Addr	1F46	8006
x"00",	-- Hex Addr	1F47	8007
x"00",	-- Hex Addr	1F48	8008
x"00",	-- Hex Addr	1F49	8009
x"00",	-- Hex Addr	1F4A	8010
x"00",	-- Hex Addr	1F4B	8011
x"00",	-- Hex Addr	1F4C	8012
x"00",	-- Hex Addr	1F4D	8013
x"00",	-- Hex Addr	1F4E	8014
x"00",	-- Hex Addr	1F4F	8015
x"00",	-- Hex Addr	1F50	8016
x"00",	-- Hex Addr	1F51	8017
x"00",	-- Hex Addr	1F52	8018
x"00",	-- Hex Addr	1F53	8019
x"00",	-- Hex Addr	1F54	8020
x"00",	-- Hex Addr	1F55	8021
x"00",	-- Hex Addr	1F56	8022
x"00",	-- Hex Addr	1F57	8023
x"00",	-- Hex Addr	1F58	8024
x"00",	-- Hex Addr	1F59	8025
x"00",	-- Hex Addr	1F5A	8026
x"00",	-- Hex Addr	1F5B	8027
x"00",	-- Hex Addr	1F5C	8028
x"00",	-- Hex Addr	1F5D	8029
x"00",	-- Hex Addr	1F5E	8030
x"00",	-- Hex Addr	1F5F	8031
x"00",	-- Hex Addr	1F60	8032
x"00",	-- Hex Addr	1F61	8033
x"00",	-- Hex Addr	1F62	8034
x"00",	-- Hex Addr	1F63	8035
x"00",	-- Hex Addr	1F64	8036
x"00",	-- Hex Addr	1F65	8037
x"00",	-- Hex Addr	1F66	8038
x"00",	-- Hex Addr	1F67	8039
x"00",	-- Hex Addr	1F68	8040
x"00",	-- Hex Addr	1F69	8041
x"00",	-- Hex Addr	1F6A	8042
x"00",	-- Hex Addr	1F6B	8043
x"00",	-- Hex Addr	1F6C	8044
x"00",	-- Hex Addr	1F6D	8045
x"00",	-- Hex Addr	1F6E	8046
x"00",	-- Hex Addr	1F6F	8047
x"00",	-- Hex Addr	1F70	8048
x"00",	-- Hex Addr	1F71	8049
x"00",	-- Hex Addr	1F72	8050
x"00",	-- Hex Addr	1F73	8051
x"00",	-- Hex Addr	1F74	8052
x"00",	-- Hex Addr	1F75	8053
x"00",	-- Hex Addr	1F76	8054
x"00",	-- Hex Addr	1F77	8055
x"00",	-- Hex Addr	1F78	8056
x"00",	-- Hex Addr	1F79	8057
x"00",	-- Hex Addr	1F7A	8058
x"00",	-- Hex Addr	1F7B	8059
x"00",	-- Hex Addr	1F7C	8060
x"00",	-- Hex Addr	1F7D	8061
x"00",	-- Hex Addr	1F7E	8062
x"00",	-- Hex Addr	1F7F	8063
x"00",	-- Hex Addr	1F80	8064
x"00",	-- Hex Addr	1F81	8065
x"00",	-- Hex Addr	1F82	8066
x"00",	-- Hex Addr	1F83	8067
x"00",	-- Hex Addr	1F84	8068
x"00",	-- Hex Addr	1F85	8069
x"00",	-- Hex Addr	1F86	8070
x"00",	-- Hex Addr	1F87	8071
x"00",	-- Hex Addr	1F88	8072
x"00",	-- Hex Addr	1F89	8073
x"00",	-- Hex Addr	1F8A	8074
x"00",	-- Hex Addr	1F8B	8075
x"00",	-- Hex Addr	1F8C	8076
x"00",	-- Hex Addr	1F8D	8077
x"00",	-- Hex Addr	1F8E	8078
x"00",	-- Hex Addr	1F8F	8079
x"00",	-- Hex Addr	1F90	8080
x"00",	-- Hex Addr	1F91	8081
x"00",	-- Hex Addr	1F92	8082
x"00",	-- Hex Addr	1F93	8083
x"00",	-- Hex Addr	1F94	8084
x"00",	-- Hex Addr	1F95	8085
x"00",	-- Hex Addr	1F96	8086
x"00",	-- Hex Addr	1F97	8087
x"00",	-- Hex Addr	1F98	8088
x"00",	-- Hex Addr	1F99	8089
x"00",	-- Hex Addr	1F9A	8090
x"00",	-- Hex Addr	1F9B	8091
x"00",	-- Hex Addr	1F9C	8092
x"00",	-- Hex Addr	1F9D	8093
x"00",	-- Hex Addr	1F9E	8094
x"00",	-- Hex Addr	1F9F	8095
x"00",	-- Hex Addr	1FA0	8096
x"00",	-- Hex Addr	1FA1	8097
x"00",	-- Hex Addr	1FA2	8098
x"00",	-- Hex Addr	1FA3	8099
x"00",	-- Hex Addr	1FA4	8100
x"00",	-- Hex Addr	1FA5	8101
x"00",	-- Hex Addr	1FA6	8102
x"00",	-- Hex Addr	1FA7	8103
x"00",	-- Hex Addr	1FA8	8104
x"00",	-- Hex Addr	1FA9	8105
x"00",	-- Hex Addr	1FAA	8106
x"00",	-- Hex Addr	1FAB	8107
x"00",	-- Hex Addr	1FAC	8108
x"00",	-- Hex Addr	1FAD	8109
x"00",	-- Hex Addr	1FAE	8110
x"00",	-- Hex Addr	1FAF	8111
x"00",	-- Hex Addr	1FB0	8112
x"00",	-- Hex Addr	1FB1	8113
x"00",	-- Hex Addr	1FB2	8114
x"00",	-- Hex Addr	1FB3	8115
x"00",	-- Hex Addr	1FB4	8116
x"00",	-- Hex Addr	1FB5	8117
x"00",	-- Hex Addr	1FB6	8118
x"00",	-- Hex Addr	1FB7	8119
x"00",	-- Hex Addr	1FB8	8120
x"00",	-- Hex Addr	1FB9	8121
x"00",	-- Hex Addr	1FBA	8122
x"00",	-- Hex Addr	1FBB	8123
x"00",	-- Hex Addr	1FBC	8124
x"00",	-- Hex Addr	1FBD	8125
x"00",	-- Hex Addr	1FBE	8126
x"00",	-- Hex Addr	1FBF	8127
x"00",	-- Hex Addr	1FC0	8128
x"00",	-- Hex Addr	1FC1	8129
x"00",	-- Hex Addr	1FC2	8130
x"00",	-- Hex Addr	1FC3	8131
x"00",	-- Hex Addr	1FC4	8132
x"00",	-- Hex Addr	1FC5	8133
x"00",	-- Hex Addr	1FC6	8134
x"00",	-- Hex Addr	1FC7	8135
x"00",	-- Hex Addr	1FC8	8136
x"00",	-- Hex Addr	1FC9	8137
x"00",	-- Hex Addr	1FCA	8138
x"00",	-- Hex Addr	1FCB	8139
x"00",	-- Hex Addr	1FCC	8140
x"00",	-- Hex Addr	1FCD	8141
x"00",	-- Hex Addr	1FCE	8142
x"00",	-- Hex Addr	1FCF	8143
x"00",	-- Hex Addr	1FD0	8144
x"00",	-- Hex Addr	1FD1	8145
x"00",	-- Hex Addr	1FD2	8146
x"00",	-- Hex Addr	1FD3	8147
x"00",	-- Hex Addr	1FD4	8148
x"00",	-- Hex Addr	1FD5	8149
x"00",	-- Hex Addr	1FD6	8150
x"00",	-- Hex Addr	1FD7	8151
x"00",	-- Hex Addr	1FD8	8152
x"00",	-- Hex Addr	1FD9	8153
x"00",	-- Hex Addr	1FDA	8154
x"00",	-- Hex Addr	1FDB	8155
x"00",	-- Hex Addr	1FDC	8156
x"00",	-- Hex Addr	1FDD	8157
x"00",	-- Hex Addr	1FDE	8158
x"00",	-- Hex Addr	1FDF	8159
x"00",	-- Hex Addr	1FE0	8160
x"00",	-- Hex Addr	1FE1	8161
x"00",	-- Hex Addr	1FE2	8162
x"00",	-- Hex Addr	1FE3	8163
x"00",	-- Hex Addr	1FE4	8164
x"00",	-- Hex Addr	1FE5	8165
x"00",	-- Hex Addr	1FE6	8166
x"00",	-- Hex Addr	1FE7	8167
x"00",	-- Hex Addr	1FE8	8168
x"00",	-- Hex Addr	1FE9	8169
x"00",	-- Hex Addr	1FEA	8170
x"00",	-- Hex Addr	1FEB	8171
x"00",	-- Hex Addr	1FEC	8172
x"00",	-- Hex Addr	1FED	8173
x"00",	-- Hex Addr	1FEE	8174
x"00",	-- Hex Addr	1FEF	8175
x"00",	-- Hex Addr	1FF0	8176
x"00",	-- Hex Addr	1FF1	8177
x"00",	-- Hex Addr	1FF2	8178
x"00",	-- Hex Addr	1FF3	8179
x"00",	-- Hex Addr	1FF4	8180
x"00",	-- Hex Addr	1FF5	8181
x"00",	-- Hex Addr	1FF6	8182
x"00",	-- Hex Addr	1FF7	8183
x"00",	-- Hex Addr	1FF8	8184
x"00",	-- Hex Addr	1FF9	8185
x"00",	-- Hex Addr	1FFA	8186
x"00",	-- Hex Addr	1FFB	8187
x"00",	-- Hex Addr	1FFC	8188
x"00",	-- Hex Addr	1FFD	8189
x"00",	-- Hex Addr	1FFE	8190
x"00",	-- Hex Addr	1FFF	8191
x"00",	-- Hex Addr	2000	8192
x"00",	-- Hex Addr	2001	8193
x"00",	-- Hex Addr	2002	8194
x"00",	-- Hex Addr	2003	8195
x"00",	-- Hex Addr	2004	8196
x"00",	-- Hex Addr	2005	8197
x"00",	-- Hex Addr	2006	8198
x"00",	-- Hex Addr	2007	8199
x"00",	-- Hex Addr	2008	8200
x"00",	-- Hex Addr	2009	8201
x"00",	-- Hex Addr	200A	8202
x"00",	-- Hex Addr	200B	8203
x"00",	-- Hex Addr	200C	8204
x"00",	-- Hex Addr	200D	8205
x"00",	-- Hex Addr	200E	8206
x"00",	-- Hex Addr	200F	8207
x"00",	-- Hex Addr	2010	8208
x"00",	-- Hex Addr	2011	8209
x"00",	-- Hex Addr	2012	8210
x"00",	-- Hex Addr	2013	8211
x"00",	-- Hex Addr	2014	8212
x"00",	-- Hex Addr	2015	8213
x"00",	-- Hex Addr	2016	8214
x"00",	-- Hex Addr	2017	8215
x"00",	-- Hex Addr	2018	8216
x"00",	-- Hex Addr	2019	8217
x"00",	-- Hex Addr	201A	8218
x"00",	-- Hex Addr	201B	8219
x"00",	-- Hex Addr	201C	8220
x"00",	-- Hex Addr	201D	8221
x"00",	-- Hex Addr	201E	8222
x"00",	-- Hex Addr	201F	8223
x"00",	-- Hex Addr	2020	8224
x"00",	-- Hex Addr	2021	8225
x"00",	-- Hex Addr	2022	8226
x"00",	-- Hex Addr	2023	8227
x"00",	-- Hex Addr	2024	8228
x"00",	-- Hex Addr	2025	8229
x"00",	-- Hex Addr	2026	8230
x"00",	-- Hex Addr	2027	8231
x"00",	-- Hex Addr	2028	8232
x"00",	-- Hex Addr	2029	8233
x"00",	-- Hex Addr	202A	8234
x"00",	-- Hex Addr	202B	8235
x"00",	-- Hex Addr	202C	8236
x"00",	-- Hex Addr	202D	8237
x"00",	-- Hex Addr	202E	8238
x"00",	-- Hex Addr	202F	8239
x"00",	-- Hex Addr	2030	8240
x"00",	-- Hex Addr	2031	8241
x"00",	-- Hex Addr	2032	8242
x"00",	-- Hex Addr	2033	8243
x"00",	-- Hex Addr	2034	8244
x"00",	-- Hex Addr	2035	8245
x"00",	-- Hex Addr	2036	8246
x"00",	-- Hex Addr	2037	8247
x"00",	-- Hex Addr	2038	8248
x"00",	-- Hex Addr	2039	8249
x"00",	-- Hex Addr	203A	8250
x"00",	-- Hex Addr	203B	8251
x"00",	-- Hex Addr	203C	8252
x"00",	-- Hex Addr	203D	8253
x"00",	-- Hex Addr	203E	8254
x"00",	-- Hex Addr	203F	8255
x"00",	-- Hex Addr	2040	8256
x"00",	-- Hex Addr	2041	8257
x"00",	-- Hex Addr	2042	8258
x"00",	-- Hex Addr	2043	8259
x"00",	-- Hex Addr	2044	8260
x"00",	-- Hex Addr	2045	8261
x"00",	-- Hex Addr	2046	8262
x"00",	-- Hex Addr	2047	8263
x"00",	-- Hex Addr	2048	8264
x"00",	-- Hex Addr	2049	8265
x"00",	-- Hex Addr	204A	8266
x"00",	-- Hex Addr	204B	8267
x"00",	-- Hex Addr	204C	8268
x"00",	-- Hex Addr	204D	8269
x"00",	-- Hex Addr	204E	8270
x"00",	-- Hex Addr	204F	8271
x"00",	-- Hex Addr	2050	8272
x"00",	-- Hex Addr	2051	8273
x"00",	-- Hex Addr	2052	8274
x"00",	-- Hex Addr	2053	8275
x"00",	-- Hex Addr	2054	8276
x"00",	-- Hex Addr	2055	8277
x"00",	-- Hex Addr	2056	8278
x"00",	-- Hex Addr	2057	8279
x"00",	-- Hex Addr	2058	8280
x"00",	-- Hex Addr	2059	8281
x"00",	-- Hex Addr	205A	8282
x"00",	-- Hex Addr	205B	8283
x"00",	-- Hex Addr	205C	8284
x"00",	-- Hex Addr	205D	8285
x"00",	-- Hex Addr	205E	8286
x"00",	-- Hex Addr	205F	8287
x"00",	-- Hex Addr	2060	8288
x"00",	-- Hex Addr	2061	8289
x"00",	-- Hex Addr	2062	8290
x"00",	-- Hex Addr	2063	8291
x"00",	-- Hex Addr	2064	8292
x"00",	-- Hex Addr	2065	8293
x"00",	-- Hex Addr	2066	8294
x"00",	-- Hex Addr	2067	8295
x"00",	-- Hex Addr	2068	8296
x"00",	-- Hex Addr	2069	8297
x"00",	-- Hex Addr	206A	8298
x"00",	-- Hex Addr	206B	8299
x"00",	-- Hex Addr	206C	8300
x"00",	-- Hex Addr	206D	8301
x"00",	-- Hex Addr	206E	8302
x"00",	-- Hex Addr	206F	8303
x"00",	-- Hex Addr	2070	8304
x"00",	-- Hex Addr	2071	8305
x"00",	-- Hex Addr	2072	8306
x"00",	-- Hex Addr	2073	8307
x"00",	-- Hex Addr	2074	8308
x"00",	-- Hex Addr	2075	8309
x"00",	-- Hex Addr	2076	8310
x"00",	-- Hex Addr	2077	8311
x"00",	-- Hex Addr	2078	8312
x"00",	-- Hex Addr	2079	8313
x"00",	-- Hex Addr	207A	8314
x"00",	-- Hex Addr	207B	8315
x"00",	-- Hex Addr	207C	8316
x"00",	-- Hex Addr	207D	8317
x"00",	-- Hex Addr	207E	8318
x"00",	-- Hex Addr	207F	8319
x"00",	-- Hex Addr	2080	8320
x"00",	-- Hex Addr	2081	8321
x"00",	-- Hex Addr	2082	8322
x"00",	-- Hex Addr	2083	8323
x"00",	-- Hex Addr	2084	8324
x"00",	-- Hex Addr	2085	8325
x"00",	-- Hex Addr	2086	8326
x"00",	-- Hex Addr	2087	8327
x"00",	-- Hex Addr	2088	8328
x"00",	-- Hex Addr	2089	8329
x"00",	-- Hex Addr	208A	8330
x"00",	-- Hex Addr	208B	8331
x"00",	-- Hex Addr	208C	8332
x"00",	-- Hex Addr	208D	8333
x"00",	-- Hex Addr	208E	8334
x"00",	-- Hex Addr	208F	8335
x"00",	-- Hex Addr	2090	8336
x"00",	-- Hex Addr	2091	8337
x"00",	-- Hex Addr	2092	8338
x"00",	-- Hex Addr	2093	8339
x"00",	-- Hex Addr	2094	8340
x"00",	-- Hex Addr	2095	8341
x"00",	-- Hex Addr	2096	8342
x"00",	-- Hex Addr	2097	8343
x"00",	-- Hex Addr	2098	8344
x"00",	-- Hex Addr	2099	8345
x"00",	-- Hex Addr	209A	8346
x"00",	-- Hex Addr	209B	8347
x"00",	-- Hex Addr	209C	8348
x"00",	-- Hex Addr	209D	8349
x"00",	-- Hex Addr	209E	8350
x"00",	-- Hex Addr	209F	8351
x"00",	-- Hex Addr	20A0	8352
x"00",	-- Hex Addr	20A1	8353
x"00",	-- Hex Addr	20A2	8354
x"00",	-- Hex Addr	20A3	8355
x"00",	-- Hex Addr	20A4	8356
x"00",	-- Hex Addr	20A5	8357
x"00",	-- Hex Addr	20A6	8358
x"00",	-- Hex Addr	20A7	8359
x"00",	-- Hex Addr	20A8	8360
x"00",	-- Hex Addr	20A9	8361
x"00",	-- Hex Addr	20AA	8362
x"00",	-- Hex Addr	20AB	8363
x"00",	-- Hex Addr	20AC	8364
x"00",	-- Hex Addr	20AD	8365
x"00",	-- Hex Addr	20AE	8366
x"00",	-- Hex Addr	20AF	8367
x"00",	-- Hex Addr	20B0	8368
x"00",	-- Hex Addr	20B1	8369
x"00",	-- Hex Addr	20B2	8370
x"00",	-- Hex Addr	20B3	8371
x"00",	-- Hex Addr	20B4	8372
x"00",	-- Hex Addr	20B5	8373
x"00",	-- Hex Addr	20B6	8374
x"00",	-- Hex Addr	20B7	8375
x"00",	-- Hex Addr	20B8	8376
x"00",	-- Hex Addr	20B9	8377
x"00",	-- Hex Addr	20BA	8378
x"00",	-- Hex Addr	20BB	8379
x"00",	-- Hex Addr	20BC	8380
x"00",	-- Hex Addr	20BD	8381
x"00",	-- Hex Addr	20BE	8382
x"00",	-- Hex Addr	20BF	8383
x"00",	-- Hex Addr	20C0	8384
x"00",	-- Hex Addr	20C1	8385
x"00",	-- Hex Addr	20C2	8386
x"00",	-- Hex Addr	20C3	8387
x"00",	-- Hex Addr	20C4	8388
x"00",	-- Hex Addr	20C5	8389
x"00",	-- Hex Addr	20C6	8390
x"00",	-- Hex Addr	20C7	8391
x"00",	-- Hex Addr	20C8	8392
x"00",	-- Hex Addr	20C9	8393
x"00",	-- Hex Addr	20CA	8394
x"00",	-- Hex Addr	20CB	8395
x"00",	-- Hex Addr	20CC	8396
x"00",	-- Hex Addr	20CD	8397
x"00",	-- Hex Addr	20CE	8398
x"00",	-- Hex Addr	20CF	8399
x"00",	-- Hex Addr	20D0	8400
x"00",	-- Hex Addr	20D1	8401
x"00",	-- Hex Addr	20D2	8402
x"00",	-- Hex Addr	20D3	8403
x"00",	-- Hex Addr	20D4	8404
x"00",	-- Hex Addr	20D5	8405
x"00",	-- Hex Addr	20D6	8406
x"00",	-- Hex Addr	20D7	8407
x"00",	-- Hex Addr	20D8	8408
x"00",	-- Hex Addr	20D9	8409
x"00",	-- Hex Addr	20DA	8410
x"00",	-- Hex Addr	20DB	8411
x"00",	-- Hex Addr	20DC	8412
x"00",	-- Hex Addr	20DD	8413
x"00",	-- Hex Addr	20DE	8414
x"00",	-- Hex Addr	20DF	8415
x"00",	-- Hex Addr	20E0	8416
x"00",	-- Hex Addr	20E1	8417
x"00",	-- Hex Addr	20E2	8418
x"00",	-- Hex Addr	20E3	8419
x"00",	-- Hex Addr	20E4	8420
x"00",	-- Hex Addr	20E5	8421
x"00",	-- Hex Addr	20E6	8422
x"00",	-- Hex Addr	20E7	8423
x"00",	-- Hex Addr	20E8	8424
x"00",	-- Hex Addr	20E9	8425
x"00",	-- Hex Addr	20EA	8426
x"00",	-- Hex Addr	20EB	8427
x"00",	-- Hex Addr	20EC	8428
x"00",	-- Hex Addr	20ED	8429
x"00",	-- Hex Addr	20EE	8430
x"00",	-- Hex Addr	20EF	8431
x"00",	-- Hex Addr	20F0	8432
x"00",	-- Hex Addr	20F1	8433
x"00",	-- Hex Addr	20F2	8434
x"00",	-- Hex Addr	20F3	8435
x"00",	-- Hex Addr	20F4	8436
x"00",	-- Hex Addr	20F5	8437
x"00",	-- Hex Addr	20F6	8438
x"00",	-- Hex Addr	20F7	8439
x"00",	-- Hex Addr	20F8	8440
x"00",	-- Hex Addr	20F9	8441
x"00",	-- Hex Addr	20FA	8442
x"00",	-- Hex Addr	20FB	8443
x"00",	-- Hex Addr	20FC	8444
x"00",	-- Hex Addr	20FD	8445
x"00",	-- Hex Addr	20FE	8446
x"00",	-- Hex Addr	20FF	8447
x"00",	-- Hex Addr	2100	8448
x"00",	-- Hex Addr	2101	8449
x"00",	-- Hex Addr	2102	8450
x"00",	-- Hex Addr	2103	8451
x"00",	-- Hex Addr	2104	8452
x"00",	-- Hex Addr	2105	8453
x"00",	-- Hex Addr	2106	8454
x"00",	-- Hex Addr	2107	8455
x"00",	-- Hex Addr	2108	8456
x"00",	-- Hex Addr	2109	8457
x"00",	-- Hex Addr	210A	8458
x"00",	-- Hex Addr	210B	8459
x"00",	-- Hex Addr	210C	8460
x"00",	-- Hex Addr	210D	8461
x"00",	-- Hex Addr	210E	8462
x"00",	-- Hex Addr	210F	8463
x"00",	-- Hex Addr	2110	8464
x"00",	-- Hex Addr	2111	8465
x"00",	-- Hex Addr	2112	8466
x"00",	-- Hex Addr	2113	8467
x"00",	-- Hex Addr	2114	8468
x"00",	-- Hex Addr	2115	8469
x"00",	-- Hex Addr	2116	8470
x"00",	-- Hex Addr	2117	8471
x"00",	-- Hex Addr	2118	8472
x"00",	-- Hex Addr	2119	8473
x"00",	-- Hex Addr	211A	8474
x"00",	-- Hex Addr	211B	8475
x"00",	-- Hex Addr	211C	8476
x"00",	-- Hex Addr	211D	8477
x"00",	-- Hex Addr	211E	8478
x"00",	-- Hex Addr	211F	8479
x"00",	-- Hex Addr	2120	8480
x"00",	-- Hex Addr	2121	8481
x"00",	-- Hex Addr	2122	8482
x"00",	-- Hex Addr	2123	8483
x"00",	-- Hex Addr	2124	8484
x"00",	-- Hex Addr	2125	8485
x"00",	-- Hex Addr	2126	8486
x"00",	-- Hex Addr	2127	8487
x"00",	-- Hex Addr	2128	8488
x"00",	-- Hex Addr	2129	8489
x"00",	-- Hex Addr	212A	8490
x"00",	-- Hex Addr	212B	8491
x"00",	-- Hex Addr	212C	8492
x"00",	-- Hex Addr	212D	8493
x"00",	-- Hex Addr	212E	8494
x"00",	-- Hex Addr	212F	8495
x"00",	-- Hex Addr	2130	8496
x"00",	-- Hex Addr	2131	8497
x"00",	-- Hex Addr	2132	8498
x"00",	-- Hex Addr	2133	8499
x"00",	-- Hex Addr	2134	8500
x"00",	-- Hex Addr	2135	8501
x"00",	-- Hex Addr	2136	8502
x"00",	-- Hex Addr	2137	8503
x"00",	-- Hex Addr	2138	8504
x"00",	-- Hex Addr	2139	8505
x"00",	-- Hex Addr	213A	8506
x"00",	-- Hex Addr	213B	8507
x"00",	-- Hex Addr	213C	8508
x"00",	-- Hex Addr	213D	8509
x"00",	-- Hex Addr	213E	8510
x"00",	-- Hex Addr	213F	8511
x"00",	-- Hex Addr	2140	8512
x"00",	-- Hex Addr	2141	8513
x"00",	-- Hex Addr	2142	8514
x"00",	-- Hex Addr	2143	8515
x"00",	-- Hex Addr	2144	8516
x"00",	-- Hex Addr	2145	8517
x"00",	-- Hex Addr	2146	8518
x"00",	-- Hex Addr	2147	8519
x"00",	-- Hex Addr	2148	8520
x"00",	-- Hex Addr	2149	8521
x"00",	-- Hex Addr	214A	8522
x"00",	-- Hex Addr	214B	8523
x"00",	-- Hex Addr	214C	8524
x"00",	-- Hex Addr	214D	8525
x"00",	-- Hex Addr	214E	8526
x"00",	-- Hex Addr	214F	8527
x"00",	-- Hex Addr	2150	8528
x"00",	-- Hex Addr	2151	8529
x"00",	-- Hex Addr	2152	8530
x"00",	-- Hex Addr	2153	8531
x"00",	-- Hex Addr	2154	8532
x"00",	-- Hex Addr	2155	8533
x"00",	-- Hex Addr	2156	8534
x"00",	-- Hex Addr	2157	8535
x"00",	-- Hex Addr	2158	8536
x"00",	-- Hex Addr	2159	8537
x"00",	-- Hex Addr	215A	8538
x"00",	-- Hex Addr	215B	8539
x"00",	-- Hex Addr	215C	8540
x"00",	-- Hex Addr	215D	8541
x"00",	-- Hex Addr	215E	8542
x"00",	-- Hex Addr	215F	8543
x"00",	-- Hex Addr	2160	8544
x"00",	-- Hex Addr	2161	8545
x"00",	-- Hex Addr	2162	8546
x"00",	-- Hex Addr	2163	8547
x"00",	-- Hex Addr	2164	8548
x"00",	-- Hex Addr	2165	8549
x"00",	-- Hex Addr	2166	8550
x"00",	-- Hex Addr	2167	8551
x"00",	-- Hex Addr	2168	8552
x"00",	-- Hex Addr	2169	8553
x"00",	-- Hex Addr	216A	8554
x"00",	-- Hex Addr	216B	8555
x"00",	-- Hex Addr	216C	8556
x"00",	-- Hex Addr	216D	8557
x"00",	-- Hex Addr	216E	8558
x"00",	-- Hex Addr	216F	8559
x"00",	-- Hex Addr	2170	8560
x"00",	-- Hex Addr	2171	8561
x"00",	-- Hex Addr	2172	8562
x"00",	-- Hex Addr	2173	8563
x"00",	-- Hex Addr	2174	8564
x"00",	-- Hex Addr	2175	8565
x"00",	-- Hex Addr	2176	8566
x"00",	-- Hex Addr	2177	8567
x"00",	-- Hex Addr	2178	8568
x"00",	-- Hex Addr	2179	8569
x"00",	-- Hex Addr	217A	8570
x"00",	-- Hex Addr	217B	8571
x"00",	-- Hex Addr	217C	8572
x"00",	-- Hex Addr	217D	8573
x"00",	-- Hex Addr	217E	8574
x"00",	-- Hex Addr	217F	8575
x"00",	-- Hex Addr	2180	8576
x"00",	-- Hex Addr	2181	8577
x"00",	-- Hex Addr	2182	8578
x"00",	-- Hex Addr	2183	8579
x"00",	-- Hex Addr	2184	8580
x"00",	-- Hex Addr	2185	8581
x"00",	-- Hex Addr	2186	8582
x"00",	-- Hex Addr	2187	8583
x"00",	-- Hex Addr	2188	8584
x"00",	-- Hex Addr	2189	8585
x"00",	-- Hex Addr	218A	8586
x"00",	-- Hex Addr	218B	8587
x"00",	-- Hex Addr	218C	8588
x"00",	-- Hex Addr	218D	8589
x"00",	-- Hex Addr	218E	8590
x"00",	-- Hex Addr	218F	8591
x"00",	-- Hex Addr	2190	8592
x"00",	-- Hex Addr	2191	8593
x"00",	-- Hex Addr	2192	8594
x"00",	-- Hex Addr	2193	8595
x"00",	-- Hex Addr	2194	8596
x"00",	-- Hex Addr	2195	8597
x"00",	-- Hex Addr	2196	8598
x"00",	-- Hex Addr	2197	8599
x"00",	-- Hex Addr	2198	8600
x"00",	-- Hex Addr	2199	8601
x"00",	-- Hex Addr	219A	8602
x"00",	-- Hex Addr	219B	8603
x"00",	-- Hex Addr	219C	8604
x"00",	-- Hex Addr	219D	8605
x"00",	-- Hex Addr	219E	8606
x"00",	-- Hex Addr	219F	8607
x"00",	-- Hex Addr	21A0	8608
x"00",	-- Hex Addr	21A1	8609
x"00",	-- Hex Addr	21A2	8610
x"00",	-- Hex Addr	21A3	8611
x"00",	-- Hex Addr	21A4	8612
x"00",	-- Hex Addr	21A5	8613
x"00",	-- Hex Addr	21A6	8614
x"00",	-- Hex Addr	21A7	8615
x"00",	-- Hex Addr	21A8	8616
x"00",	-- Hex Addr	21A9	8617
x"00",	-- Hex Addr	21AA	8618
x"00",	-- Hex Addr	21AB	8619
x"00",	-- Hex Addr	21AC	8620
x"00",	-- Hex Addr	21AD	8621
x"00",	-- Hex Addr	21AE	8622
x"00",	-- Hex Addr	21AF	8623
x"00",	-- Hex Addr	21B0	8624
x"00",	-- Hex Addr	21B1	8625
x"00",	-- Hex Addr	21B2	8626
x"00",	-- Hex Addr	21B3	8627
x"00",	-- Hex Addr	21B4	8628
x"00",	-- Hex Addr	21B5	8629
x"00",	-- Hex Addr	21B6	8630
x"00",	-- Hex Addr	21B7	8631
x"00",	-- Hex Addr	21B8	8632
x"00",	-- Hex Addr	21B9	8633
x"00",	-- Hex Addr	21BA	8634
x"00",	-- Hex Addr	21BB	8635
x"00",	-- Hex Addr	21BC	8636
x"00",	-- Hex Addr	21BD	8637
x"00",	-- Hex Addr	21BE	8638
x"00",	-- Hex Addr	21BF	8639
x"00",	-- Hex Addr	21C0	8640
x"00",	-- Hex Addr	21C1	8641
x"00",	-- Hex Addr	21C2	8642
x"00",	-- Hex Addr	21C3	8643
x"00",	-- Hex Addr	21C4	8644
x"00",	-- Hex Addr	21C5	8645
x"00",	-- Hex Addr	21C6	8646
x"00",	-- Hex Addr	21C7	8647
x"00",	-- Hex Addr	21C8	8648
x"00",	-- Hex Addr	21C9	8649
x"00",	-- Hex Addr	21CA	8650
x"00",	-- Hex Addr	21CB	8651
x"00",	-- Hex Addr	21CC	8652
x"00",	-- Hex Addr	21CD	8653
x"00",	-- Hex Addr	21CE	8654
x"00",	-- Hex Addr	21CF	8655
x"00",	-- Hex Addr	21D0	8656
x"00",	-- Hex Addr	21D1	8657
x"00",	-- Hex Addr	21D2	8658
x"00",	-- Hex Addr	21D3	8659
x"00",	-- Hex Addr	21D4	8660
x"00",	-- Hex Addr	21D5	8661
x"00",	-- Hex Addr	21D6	8662
x"00",	-- Hex Addr	21D7	8663
x"00",	-- Hex Addr	21D8	8664
x"00",	-- Hex Addr	21D9	8665
x"00",	-- Hex Addr	21DA	8666
x"00",	-- Hex Addr	21DB	8667
x"00",	-- Hex Addr	21DC	8668
x"00",	-- Hex Addr	21DD	8669
x"00",	-- Hex Addr	21DE	8670
x"00",	-- Hex Addr	21DF	8671
x"00",	-- Hex Addr	21E0	8672
x"00",	-- Hex Addr	21E1	8673
x"00",	-- Hex Addr	21E2	8674
x"00",	-- Hex Addr	21E3	8675
x"00",	-- Hex Addr	21E4	8676
x"00",	-- Hex Addr	21E5	8677
x"00",	-- Hex Addr	21E6	8678
x"00",	-- Hex Addr	21E7	8679
x"00",	-- Hex Addr	21E8	8680
x"00",	-- Hex Addr	21E9	8681
x"00",	-- Hex Addr	21EA	8682
x"00",	-- Hex Addr	21EB	8683
x"00",	-- Hex Addr	21EC	8684
x"00",	-- Hex Addr	21ED	8685
x"00",	-- Hex Addr	21EE	8686
x"00",	-- Hex Addr	21EF	8687
x"00",	-- Hex Addr	21F0	8688
x"00",	-- Hex Addr	21F1	8689
x"00",	-- Hex Addr	21F2	8690
x"00",	-- Hex Addr	21F3	8691
x"00",	-- Hex Addr	21F4	8692
x"00",	-- Hex Addr	21F5	8693
x"00",	-- Hex Addr	21F6	8694
x"00",	-- Hex Addr	21F7	8695
x"00",	-- Hex Addr	21F8	8696
x"00",	-- Hex Addr	21F9	8697
x"00",	-- Hex Addr	21FA	8698
x"00",	-- Hex Addr	21FB	8699
x"00",	-- Hex Addr	21FC	8700
x"00",	-- Hex Addr	21FD	8701
x"00",	-- Hex Addr	21FE	8702
x"00",	-- Hex Addr	21FF	8703
x"00",	-- Hex Addr	2200	8704
x"00",	-- Hex Addr	2201	8705
x"00",	-- Hex Addr	2202	8706
x"00",	-- Hex Addr	2203	8707
x"00",	-- Hex Addr	2204	8708
x"00",	-- Hex Addr	2205	8709
x"00",	-- Hex Addr	2206	8710
x"00",	-- Hex Addr	2207	8711
x"00",	-- Hex Addr	2208	8712
x"00",	-- Hex Addr	2209	8713
x"00",	-- Hex Addr	220A	8714
x"00",	-- Hex Addr	220B	8715
x"00",	-- Hex Addr	220C	8716
x"00",	-- Hex Addr	220D	8717
x"00",	-- Hex Addr	220E	8718
x"00",	-- Hex Addr	220F	8719
x"00",	-- Hex Addr	2210	8720
x"00",	-- Hex Addr	2211	8721
x"00",	-- Hex Addr	2212	8722
x"00",	-- Hex Addr	2213	8723
x"00",	-- Hex Addr	2214	8724
x"00",	-- Hex Addr	2215	8725
x"00",	-- Hex Addr	2216	8726
x"00",	-- Hex Addr	2217	8727
x"00",	-- Hex Addr	2218	8728
x"00",	-- Hex Addr	2219	8729
x"00",	-- Hex Addr	221A	8730
x"00",	-- Hex Addr	221B	8731
x"00",	-- Hex Addr	221C	8732
x"00",	-- Hex Addr	221D	8733
x"00",	-- Hex Addr	221E	8734
x"00",	-- Hex Addr	221F	8735
x"00",	-- Hex Addr	2220	8736
x"00",	-- Hex Addr	2221	8737
x"00",	-- Hex Addr	2222	8738
x"00",	-- Hex Addr	2223	8739
x"00",	-- Hex Addr	2224	8740
x"00",	-- Hex Addr	2225	8741
x"00",	-- Hex Addr	2226	8742
x"00",	-- Hex Addr	2227	8743
x"00",	-- Hex Addr	2228	8744
x"00",	-- Hex Addr	2229	8745
x"00",	-- Hex Addr	222A	8746
x"00",	-- Hex Addr	222B	8747
x"00",	-- Hex Addr	222C	8748
x"00",	-- Hex Addr	222D	8749
x"00",	-- Hex Addr	222E	8750
x"00",	-- Hex Addr	222F	8751
x"00",	-- Hex Addr	2230	8752
x"00",	-- Hex Addr	2231	8753
x"00",	-- Hex Addr	2232	8754
x"00",	-- Hex Addr	2233	8755
x"00",	-- Hex Addr	2234	8756
x"00",	-- Hex Addr	2235	8757
x"00",	-- Hex Addr	2236	8758
x"00",	-- Hex Addr	2237	8759
x"00",	-- Hex Addr	2238	8760
x"00",	-- Hex Addr	2239	8761
x"00",	-- Hex Addr	223A	8762
x"00",	-- Hex Addr	223B	8763
x"00",	-- Hex Addr	223C	8764
x"00",	-- Hex Addr	223D	8765
x"00",	-- Hex Addr	223E	8766
x"00",	-- Hex Addr	223F	8767
x"00",	-- Hex Addr	2240	8768
x"00",	-- Hex Addr	2241	8769
x"00",	-- Hex Addr	2242	8770
x"00",	-- Hex Addr	2243	8771
x"00",	-- Hex Addr	2244	8772
x"00",	-- Hex Addr	2245	8773
x"00",	-- Hex Addr	2246	8774
x"00",	-- Hex Addr	2247	8775
x"00",	-- Hex Addr	2248	8776
x"00",	-- Hex Addr	2249	8777
x"00",	-- Hex Addr	224A	8778
x"00",	-- Hex Addr	224B	8779
x"00",	-- Hex Addr	224C	8780
x"00",	-- Hex Addr	224D	8781
x"00",	-- Hex Addr	224E	8782
x"00",	-- Hex Addr	224F	8783
x"00",	-- Hex Addr	2250	8784
x"00",	-- Hex Addr	2251	8785
x"00",	-- Hex Addr	2252	8786
x"00",	-- Hex Addr	2253	8787
x"00",	-- Hex Addr	2254	8788
x"00",	-- Hex Addr	2255	8789
x"00",	-- Hex Addr	2256	8790
x"00",	-- Hex Addr	2257	8791
x"00",	-- Hex Addr	2258	8792
x"00",	-- Hex Addr	2259	8793
x"00",	-- Hex Addr	225A	8794
x"00",	-- Hex Addr	225B	8795
x"00",	-- Hex Addr	225C	8796
x"00",	-- Hex Addr	225D	8797
x"00",	-- Hex Addr	225E	8798
x"00",	-- Hex Addr	225F	8799
x"00",	-- Hex Addr	2260	8800
x"00",	-- Hex Addr	2261	8801
x"00",	-- Hex Addr	2262	8802
x"00",	-- Hex Addr	2263	8803
x"00",	-- Hex Addr	2264	8804
x"00",	-- Hex Addr	2265	8805
x"00",	-- Hex Addr	2266	8806
x"00",	-- Hex Addr	2267	8807
x"00",	-- Hex Addr	2268	8808
x"00",	-- Hex Addr	2269	8809
x"00",	-- Hex Addr	226A	8810
x"00",	-- Hex Addr	226B	8811
x"00",	-- Hex Addr	226C	8812
x"00",	-- Hex Addr	226D	8813
x"00",	-- Hex Addr	226E	8814
x"00",	-- Hex Addr	226F	8815
x"00",	-- Hex Addr	2270	8816
x"00",	-- Hex Addr	2271	8817
x"00",	-- Hex Addr	2272	8818
x"00",	-- Hex Addr	2273	8819
x"00",	-- Hex Addr	2274	8820
x"00",	-- Hex Addr	2275	8821
x"00",	-- Hex Addr	2276	8822
x"00",	-- Hex Addr	2277	8823
x"00",	-- Hex Addr	2278	8824
x"00",	-- Hex Addr	2279	8825
x"00",	-- Hex Addr	227A	8826
x"00",	-- Hex Addr	227B	8827
x"00",	-- Hex Addr	227C	8828
x"00",	-- Hex Addr	227D	8829
x"00",	-- Hex Addr	227E	8830
x"00",	-- Hex Addr	227F	8831
x"00",	-- Hex Addr	2280	8832
x"00",	-- Hex Addr	2281	8833
x"00",	-- Hex Addr	2282	8834
x"00",	-- Hex Addr	2283	8835
x"00",	-- Hex Addr	2284	8836
x"00",	-- Hex Addr	2285	8837
x"00",	-- Hex Addr	2286	8838
x"00",	-- Hex Addr	2287	8839
x"00",	-- Hex Addr	2288	8840
x"00",	-- Hex Addr	2289	8841
x"00",	-- Hex Addr	228A	8842
x"00",	-- Hex Addr	228B	8843
x"00",	-- Hex Addr	228C	8844
x"00",	-- Hex Addr	228D	8845
x"00",	-- Hex Addr	228E	8846
x"00",	-- Hex Addr	228F	8847
x"00",	-- Hex Addr	2290	8848
x"00",	-- Hex Addr	2291	8849
x"00",	-- Hex Addr	2292	8850
x"00",	-- Hex Addr	2293	8851
x"00",	-- Hex Addr	2294	8852
x"00",	-- Hex Addr	2295	8853
x"00",	-- Hex Addr	2296	8854
x"00",	-- Hex Addr	2297	8855
x"00",	-- Hex Addr	2298	8856
x"00",	-- Hex Addr	2299	8857
x"00",	-- Hex Addr	229A	8858
x"00",	-- Hex Addr	229B	8859
x"00",	-- Hex Addr	229C	8860
x"00",	-- Hex Addr	229D	8861
x"00",	-- Hex Addr	229E	8862
x"00",	-- Hex Addr	229F	8863
x"00",	-- Hex Addr	22A0	8864
x"00",	-- Hex Addr	22A1	8865
x"00",	-- Hex Addr	22A2	8866
x"00",	-- Hex Addr	22A3	8867
x"00",	-- Hex Addr	22A4	8868
x"00",	-- Hex Addr	22A5	8869
x"00",	-- Hex Addr	22A6	8870
x"00",	-- Hex Addr	22A7	8871
x"00",	-- Hex Addr	22A8	8872
x"00",	-- Hex Addr	22A9	8873
x"00",	-- Hex Addr	22AA	8874
x"00",	-- Hex Addr	22AB	8875
x"00",	-- Hex Addr	22AC	8876
x"00",	-- Hex Addr	22AD	8877
x"00",	-- Hex Addr	22AE	8878
x"00",	-- Hex Addr	22AF	8879
x"00",	-- Hex Addr	22B0	8880
x"00",	-- Hex Addr	22B1	8881
x"00",	-- Hex Addr	22B2	8882
x"00",	-- Hex Addr	22B3	8883
x"00",	-- Hex Addr	22B4	8884
x"00",	-- Hex Addr	22B5	8885
x"00",	-- Hex Addr	22B6	8886
x"00",	-- Hex Addr	22B7	8887
x"00",	-- Hex Addr	22B8	8888
x"00",	-- Hex Addr	22B9	8889
x"00",	-- Hex Addr	22BA	8890
x"00",	-- Hex Addr	22BB	8891
x"00",	-- Hex Addr	22BC	8892
x"00",	-- Hex Addr	22BD	8893
x"00",	-- Hex Addr	22BE	8894
x"00",	-- Hex Addr	22BF	8895
x"00",	-- Hex Addr	22C0	8896
x"00",	-- Hex Addr	22C1	8897
x"00",	-- Hex Addr	22C2	8898
x"00",	-- Hex Addr	22C3	8899
x"00",	-- Hex Addr	22C4	8900
x"00",	-- Hex Addr	22C5	8901
x"00",	-- Hex Addr	22C6	8902
x"00",	-- Hex Addr	22C7	8903
x"00",	-- Hex Addr	22C8	8904
x"00",	-- Hex Addr	22C9	8905
x"00",	-- Hex Addr	22CA	8906
x"00",	-- Hex Addr	22CB	8907
x"00",	-- Hex Addr	22CC	8908
x"00",	-- Hex Addr	22CD	8909
x"00",	-- Hex Addr	22CE	8910
x"00",	-- Hex Addr	22CF	8911
x"00",	-- Hex Addr	22D0	8912
x"00",	-- Hex Addr	22D1	8913
x"00",	-- Hex Addr	22D2	8914
x"00",	-- Hex Addr	22D3	8915
x"00",	-- Hex Addr	22D4	8916
x"00",	-- Hex Addr	22D5	8917
x"00",	-- Hex Addr	22D6	8918
x"00",	-- Hex Addr	22D7	8919
x"00",	-- Hex Addr	22D8	8920
x"00",	-- Hex Addr	22D9	8921
x"00",	-- Hex Addr	22DA	8922
x"00",	-- Hex Addr	22DB	8923
x"00",	-- Hex Addr	22DC	8924
x"00",	-- Hex Addr	22DD	8925
x"00",	-- Hex Addr	22DE	8926
x"00",	-- Hex Addr	22DF	8927
x"00",	-- Hex Addr	22E0	8928
x"00",	-- Hex Addr	22E1	8929
x"00",	-- Hex Addr	22E2	8930
x"00",	-- Hex Addr	22E3	8931
x"00",	-- Hex Addr	22E4	8932
x"00",	-- Hex Addr	22E5	8933
x"00",	-- Hex Addr	22E6	8934
x"00",	-- Hex Addr	22E7	8935
x"00",	-- Hex Addr	22E8	8936
x"00",	-- Hex Addr	22E9	8937
x"00",	-- Hex Addr	22EA	8938
x"00",	-- Hex Addr	22EB	8939
x"00",	-- Hex Addr	22EC	8940
x"00",	-- Hex Addr	22ED	8941
x"00",	-- Hex Addr	22EE	8942
x"00",	-- Hex Addr	22EF	8943
x"00",	-- Hex Addr	22F0	8944
x"00",	-- Hex Addr	22F1	8945
x"00",	-- Hex Addr	22F2	8946
x"00",	-- Hex Addr	22F3	8947
x"00",	-- Hex Addr	22F4	8948
x"00",	-- Hex Addr	22F5	8949
x"00",	-- Hex Addr	22F6	8950
x"00",	-- Hex Addr	22F7	8951
x"00",	-- Hex Addr	22F8	8952
x"00",	-- Hex Addr	22F9	8953
x"00",	-- Hex Addr	22FA	8954
x"00",	-- Hex Addr	22FB	8955
x"00",	-- Hex Addr	22FC	8956
x"00",	-- Hex Addr	22FD	8957
x"00",	-- Hex Addr	22FE	8958
x"00",	-- Hex Addr	22FF	8959
x"00",	-- Hex Addr	2300	8960
x"00",	-- Hex Addr	2301	8961
x"00",	-- Hex Addr	2302	8962
x"00",	-- Hex Addr	2303	8963
x"00",	-- Hex Addr	2304	8964
x"00",	-- Hex Addr	2305	8965
x"00",	-- Hex Addr	2306	8966
x"00",	-- Hex Addr	2307	8967
x"00",	-- Hex Addr	2308	8968
x"00",	-- Hex Addr	2309	8969
x"00",	-- Hex Addr	230A	8970
x"00",	-- Hex Addr	230B	8971
x"00",	-- Hex Addr	230C	8972
x"00",	-- Hex Addr	230D	8973
x"00",	-- Hex Addr	230E	8974
x"00",	-- Hex Addr	230F	8975
x"00",	-- Hex Addr	2310	8976
x"00",	-- Hex Addr	2311	8977
x"00",	-- Hex Addr	2312	8978
x"00",	-- Hex Addr	2313	8979
x"00",	-- Hex Addr	2314	8980
x"00",	-- Hex Addr	2315	8981
x"00",	-- Hex Addr	2316	8982
x"00",	-- Hex Addr	2317	8983
x"00",	-- Hex Addr	2318	8984
x"00",	-- Hex Addr	2319	8985
x"00",	-- Hex Addr	231A	8986
x"00",	-- Hex Addr	231B	8987
x"00",	-- Hex Addr	231C	8988
x"00",	-- Hex Addr	231D	8989
x"00",	-- Hex Addr	231E	8990
x"00",	-- Hex Addr	231F	8991
x"00",	-- Hex Addr	2320	8992
x"00",	-- Hex Addr	2321	8993
x"00",	-- Hex Addr	2322	8994
x"00",	-- Hex Addr	2323	8995
x"00",	-- Hex Addr	2324	8996
x"00",	-- Hex Addr	2325	8997
x"00",	-- Hex Addr	2326	8998
x"00",	-- Hex Addr	2327	8999
x"00",	-- Hex Addr	2328	9000
x"00",	-- Hex Addr	2329	9001
x"00",	-- Hex Addr	232A	9002
x"00",	-- Hex Addr	232B	9003
x"00",	-- Hex Addr	232C	9004
x"00",	-- Hex Addr	232D	9005
x"00",	-- Hex Addr	232E	9006
x"00",	-- Hex Addr	232F	9007
x"00",	-- Hex Addr	2330	9008
x"00",	-- Hex Addr	2331	9009
x"00",	-- Hex Addr	2332	9010
x"00",	-- Hex Addr	2333	9011
x"00",	-- Hex Addr	2334	9012
x"00",	-- Hex Addr	2335	9013
x"00",	-- Hex Addr	2336	9014
x"00",	-- Hex Addr	2337	9015
x"00",	-- Hex Addr	2338	9016
x"00",	-- Hex Addr	2339	9017
x"00",	-- Hex Addr	233A	9018
x"00",	-- Hex Addr	233B	9019
x"00",	-- Hex Addr	233C	9020
x"00",	-- Hex Addr	233D	9021
x"00",	-- Hex Addr	233E	9022
x"00",	-- Hex Addr	233F	9023
x"00",	-- Hex Addr	2340	9024
x"00",	-- Hex Addr	2341	9025
x"00",	-- Hex Addr	2342	9026
x"00",	-- Hex Addr	2343	9027
x"00",	-- Hex Addr	2344	9028
x"00",	-- Hex Addr	2345	9029
x"00",	-- Hex Addr	2346	9030
x"00",	-- Hex Addr	2347	9031
x"00",	-- Hex Addr	2348	9032
x"00",	-- Hex Addr	2349	9033
x"00",	-- Hex Addr	234A	9034
x"00",	-- Hex Addr	234B	9035
x"00",	-- Hex Addr	234C	9036
x"00",	-- Hex Addr	234D	9037
x"00",	-- Hex Addr	234E	9038
x"00",	-- Hex Addr	234F	9039
x"00",	-- Hex Addr	2350	9040
x"00",	-- Hex Addr	2351	9041
x"00",	-- Hex Addr	2352	9042
x"00",	-- Hex Addr	2353	9043
x"00",	-- Hex Addr	2354	9044
x"00",	-- Hex Addr	2355	9045
x"00",	-- Hex Addr	2356	9046
x"00",	-- Hex Addr	2357	9047
x"00",	-- Hex Addr	2358	9048
x"00",	-- Hex Addr	2359	9049
x"00",	-- Hex Addr	235A	9050
x"00",	-- Hex Addr	235B	9051
x"00",	-- Hex Addr	235C	9052
x"00",	-- Hex Addr	235D	9053
x"00",	-- Hex Addr	235E	9054
x"00",	-- Hex Addr	235F	9055
x"00",	-- Hex Addr	2360	9056
x"00",	-- Hex Addr	2361	9057
x"00",	-- Hex Addr	2362	9058
x"00",	-- Hex Addr	2363	9059
x"00",	-- Hex Addr	2364	9060
x"00",	-- Hex Addr	2365	9061
x"00",	-- Hex Addr	2366	9062
x"00",	-- Hex Addr	2367	9063
x"00",	-- Hex Addr	2368	9064
x"00",	-- Hex Addr	2369	9065
x"00",	-- Hex Addr	236A	9066
x"00",	-- Hex Addr	236B	9067
x"00",	-- Hex Addr	236C	9068
x"00",	-- Hex Addr	236D	9069
x"00",	-- Hex Addr	236E	9070
x"00",	-- Hex Addr	236F	9071
x"00",	-- Hex Addr	2370	9072
x"00",	-- Hex Addr	2371	9073
x"00",	-- Hex Addr	2372	9074
x"00",	-- Hex Addr	2373	9075
x"00",	-- Hex Addr	2374	9076
x"00",	-- Hex Addr	2375	9077
x"00",	-- Hex Addr	2376	9078
x"00",	-- Hex Addr	2377	9079
x"00",	-- Hex Addr	2378	9080
x"00",	-- Hex Addr	2379	9081
x"00",	-- Hex Addr	237A	9082
x"00",	-- Hex Addr	237B	9083
x"00",	-- Hex Addr	237C	9084
x"00",	-- Hex Addr	237D	9085
x"00",	-- Hex Addr	237E	9086
x"00",	-- Hex Addr	237F	9087
x"00",	-- Hex Addr	2380	9088
x"00",	-- Hex Addr	2381	9089
x"00",	-- Hex Addr	2382	9090
x"00",	-- Hex Addr	2383	9091
x"00",	-- Hex Addr	2384	9092
x"00",	-- Hex Addr	2385	9093
x"00",	-- Hex Addr	2386	9094
x"00",	-- Hex Addr	2387	9095
x"00",	-- Hex Addr	2388	9096
x"00",	-- Hex Addr	2389	9097
x"00",	-- Hex Addr	238A	9098
x"00",	-- Hex Addr	238B	9099
x"00",	-- Hex Addr	238C	9100
x"00",	-- Hex Addr	238D	9101
x"00",	-- Hex Addr	238E	9102
x"00",	-- Hex Addr	238F	9103
x"00",	-- Hex Addr	2390	9104
x"00",	-- Hex Addr	2391	9105
x"00",	-- Hex Addr	2392	9106
x"00",	-- Hex Addr	2393	9107
x"00",	-- Hex Addr	2394	9108
x"00",	-- Hex Addr	2395	9109
x"00",	-- Hex Addr	2396	9110
x"00",	-- Hex Addr	2397	9111
x"00",	-- Hex Addr	2398	9112
x"00",	-- Hex Addr	2399	9113
x"00",	-- Hex Addr	239A	9114
x"00",	-- Hex Addr	239B	9115
x"00",	-- Hex Addr	239C	9116
x"00",	-- Hex Addr	239D	9117
x"00",	-- Hex Addr	239E	9118
x"00",	-- Hex Addr	239F	9119
x"00",	-- Hex Addr	23A0	9120
x"00",	-- Hex Addr	23A1	9121
x"00",	-- Hex Addr	23A2	9122
x"00",	-- Hex Addr	23A3	9123
x"00",	-- Hex Addr	23A4	9124
x"00",	-- Hex Addr	23A5	9125
x"00",	-- Hex Addr	23A6	9126
x"00",	-- Hex Addr	23A7	9127
x"00",	-- Hex Addr	23A8	9128
x"00",	-- Hex Addr	23A9	9129
x"00",	-- Hex Addr	23AA	9130
x"00",	-- Hex Addr	23AB	9131
x"00",	-- Hex Addr	23AC	9132
x"00",	-- Hex Addr	23AD	9133
x"00",	-- Hex Addr	23AE	9134
x"00",	-- Hex Addr	23AF	9135
x"00",	-- Hex Addr	23B0	9136
x"00",	-- Hex Addr	23B1	9137
x"00",	-- Hex Addr	23B2	9138
x"00",	-- Hex Addr	23B3	9139
x"00",	-- Hex Addr	23B4	9140
x"00",	-- Hex Addr	23B5	9141
x"00",	-- Hex Addr	23B6	9142
x"00",	-- Hex Addr	23B7	9143
x"00",	-- Hex Addr	23B8	9144
x"00",	-- Hex Addr	23B9	9145
x"00",	-- Hex Addr	23BA	9146
x"00",	-- Hex Addr	23BB	9147
x"00",	-- Hex Addr	23BC	9148
x"00",	-- Hex Addr	23BD	9149
x"00",	-- Hex Addr	23BE	9150
x"00",	-- Hex Addr	23BF	9151
x"00",	-- Hex Addr	23C0	9152
x"00",	-- Hex Addr	23C1	9153
x"00",	-- Hex Addr	23C2	9154
x"00",	-- Hex Addr	23C3	9155
x"00",	-- Hex Addr	23C4	9156
x"00",	-- Hex Addr	23C5	9157
x"00",	-- Hex Addr	23C6	9158
x"00",	-- Hex Addr	23C7	9159
x"00",	-- Hex Addr	23C8	9160
x"00",	-- Hex Addr	23C9	9161
x"00",	-- Hex Addr	23CA	9162
x"00",	-- Hex Addr	23CB	9163
x"00",	-- Hex Addr	23CC	9164
x"00",	-- Hex Addr	23CD	9165
x"00",	-- Hex Addr	23CE	9166
x"00",	-- Hex Addr	23CF	9167
x"00",	-- Hex Addr	23D0	9168
x"00",	-- Hex Addr	23D1	9169
x"00",	-- Hex Addr	23D2	9170
x"00",	-- Hex Addr	23D3	9171
x"00",	-- Hex Addr	23D4	9172
x"00",	-- Hex Addr	23D5	9173
x"00",	-- Hex Addr	23D6	9174
x"00",	-- Hex Addr	23D7	9175
x"00",	-- Hex Addr	23D8	9176
x"00",	-- Hex Addr	23D9	9177
x"00",	-- Hex Addr	23DA	9178
x"00",	-- Hex Addr	23DB	9179
x"00",	-- Hex Addr	23DC	9180
x"00",	-- Hex Addr	23DD	9181
x"00",	-- Hex Addr	23DE	9182
x"00",	-- Hex Addr	23DF	9183
x"00",	-- Hex Addr	23E0	9184
x"00",	-- Hex Addr	23E1	9185
x"00",	-- Hex Addr	23E2	9186
x"00",	-- Hex Addr	23E3	9187
x"00",	-- Hex Addr	23E4	9188
x"00",	-- Hex Addr	23E5	9189
x"00",	-- Hex Addr	23E6	9190
x"00",	-- Hex Addr	23E7	9191
x"00",	-- Hex Addr	23E8	9192
x"00",	-- Hex Addr	23E9	9193
x"00",	-- Hex Addr	23EA	9194
x"00",	-- Hex Addr	23EB	9195
x"00",	-- Hex Addr	23EC	9196
x"00",	-- Hex Addr	23ED	9197
x"00",	-- Hex Addr	23EE	9198
x"00",	-- Hex Addr	23EF	9199
x"00",	-- Hex Addr	23F0	9200
x"00",	-- Hex Addr	23F1	9201
x"00",	-- Hex Addr	23F2	9202
x"00",	-- Hex Addr	23F3	9203
x"00",	-- Hex Addr	23F4	9204
x"00",	-- Hex Addr	23F5	9205
x"00",	-- Hex Addr	23F6	9206
x"00",	-- Hex Addr	23F7	9207
x"00",	-- Hex Addr	23F8	9208
x"00",	-- Hex Addr	23F9	9209
x"00",	-- Hex Addr	23FA	9210
x"00",	-- Hex Addr	23FB	9211
x"00",	-- Hex Addr	23FC	9212
x"00",	-- Hex Addr	23FD	9213
x"00",	-- Hex Addr	23FE	9214
x"00",	-- Hex Addr	23FF	9215
x"00",	-- Hex Addr	2400	9216
x"00",	-- Hex Addr	2401	9217
x"00",	-- Hex Addr	2402	9218
x"00",	-- Hex Addr	2403	9219
x"00",	-- Hex Addr	2404	9220
x"00",	-- Hex Addr	2405	9221
x"00",	-- Hex Addr	2406	9222
x"00",	-- Hex Addr	2407	9223
x"00",	-- Hex Addr	2408	9224
x"00",	-- Hex Addr	2409	9225
x"00",	-- Hex Addr	240A	9226
x"00",	-- Hex Addr	240B	9227
x"00",	-- Hex Addr	240C	9228
x"00",	-- Hex Addr	240D	9229
x"00",	-- Hex Addr	240E	9230
x"00",	-- Hex Addr	240F	9231
x"00",	-- Hex Addr	2410	9232
x"00",	-- Hex Addr	2411	9233
x"00",	-- Hex Addr	2412	9234
x"00",	-- Hex Addr	2413	9235
x"00",	-- Hex Addr	2414	9236
x"00",	-- Hex Addr	2415	9237
x"00",	-- Hex Addr	2416	9238
x"00",	-- Hex Addr	2417	9239
x"00",	-- Hex Addr	2418	9240
x"00",	-- Hex Addr	2419	9241
x"00",	-- Hex Addr	241A	9242
x"00",	-- Hex Addr	241B	9243
x"00",	-- Hex Addr	241C	9244
x"00",	-- Hex Addr	241D	9245
x"00",	-- Hex Addr	241E	9246
x"00",	-- Hex Addr	241F	9247
x"00",	-- Hex Addr	2420	9248
x"00",	-- Hex Addr	2421	9249
x"00",	-- Hex Addr	2422	9250
x"00",	-- Hex Addr	2423	9251
x"00",	-- Hex Addr	2424	9252
x"00",	-- Hex Addr	2425	9253
x"00",	-- Hex Addr	2426	9254
x"00",	-- Hex Addr	2427	9255
x"00",	-- Hex Addr	2428	9256
x"00",	-- Hex Addr	2429	9257
x"00",	-- Hex Addr	242A	9258
x"00",	-- Hex Addr	242B	9259
x"00",	-- Hex Addr	242C	9260
x"00",	-- Hex Addr	242D	9261
x"00",	-- Hex Addr	242E	9262
x"00",	-- Hex Addr	242F	9263
x"00",	-- Hex Addr	2430	9264
x"00",	-- Hex Addr	2431	9265
x"00",	-- Hex Addr	2432	9266
x"00",	-- Hex Addr	2433	9267
x"00",	-- Hex Addr	2434	9268
x"00",	-- Hex Addr	2435	9269
x"00",	-- Hex Addr	2436	9270
x"00",	-- Hex Addr	2437	9271
x"00",	-- Hex Addr	2438	9272
x"00",	-- Hex Addr	2439	9273
x"00",	-- Hex Addr	243A	9274
x"00",	-- Hex Addr	243B	9275
x"00",	-- Hex Addr	243C	9276
x"00",	-- Hex Addr	243D	9277
x"00",	-- Hex Addr	243E	9278
x"00",	-- Hex Addr	243F	9279
x"00",	-- Hex Addr	2440	9280
x"00",	-- Hex Addr	2441	9281
x"00",	-- Hex Addr	2442	9282
x"00",	-- Hex Addr	2443	9283
x"00",	-- Hex Addr	2444	9284
x"00",	-- Hex Addr	2445	9285
x"00",	-- Hex Addr	2446	9286
x"00",	-- Hex Addr	2447	9287
x"00",	-- Hex Addr	2448	9288
x"00",	-- Hex Addr	2449	9289
x"00",	-- Hex Addr	244A	9290
x"00",	-- Hex Addr	244B	9291
x"00",	-- Hex Addr	244C	9292
x"00",	-- Hex Addr	244D	9293
x"00",	-- Hex Addr	244E	9294
x"00",	-- Hex Addr	244F	9295
x"00",	-- Hex Addr	2450	9296
x"00",	-- Hex Addr	2451	9297
x"00",	-- Hex Addr	2452	9298
x"00",	-- Hex Addr	2453	9299
x"00",	-- Hex Addr	2454	9300
x"00",	-- Hex Addr	2455	9301
x"00",	-- Hex Addr	2456	9302
x"00",	-- Hex Addr	2457	9303
x"00",	-- Hex Addr	2458	9304
x"00",	-- Hex Addr	2459	9305
x"00",	-- Hex Addr	245A	9306
x"00",	-- Hex Addr	245B	9307
x"00",	-- Hex Addr	245C	9308
x"00",	-- Hex Addr	245D	9309
x"00",	-- Hex Addr	245E	9310
x"00",	-- Hex Addr	245F	9311
x"00",	-- Hex Addr	2460	9312
x"00",	-- Hex Addr	2461	9313
x"00",	-- Hex Addr	2462	9314
x"00",	-- Hex Addr	2463	9315
x"00",	-- Hex Addr	2464	9316
x"00",	-- Hex Addr	2465	9317
x"00",	-- Hex Addr	2466	9318
x"00",	-- Hex Addr	2467	9319
x"00",	-- Hex Addr	2468	9320
x"00",	-- Hex Addr	2469	9321
x"00",	-- Hex Addr	246A	9322
x"00",	-- Hex Addr	246B	9323
x"00",	-- Hex Addr	246C	9324
x"00",	-- Hex Addr	246D	9325
x"00",	-- Hex Addr	246E	9326
x"00",	-- Hex Addr	246F	9327
x"00",	-- Hex Addr	2470	9328
x"00",	-- Hex Addr	2471	9329
x"00",	-- Hex Addr	2472	9330
x"00",	-- Hex Addr	2473	9331
x"00",	-- Hex Addr	2474	9332
x"00",	-- Hex Addr	2475	9333
x"00",	-- Hex Addr	2476	9334
x"00",	-- Hex Addr	2477	9335
x"00",	-- Hex Addr	2478	9336
x"00",	-- Hex Addr	2479	9337
x"00",	-- Hex Addr	247A	9338
x"00",	-- Hex Addr	247B	9339
x"00",	-- Hex Addr	247C	9340
x"00",	-- Hex Addr	247D	9341
x"00",	-- Hex Addr	247E	9342
x"00",	-- Hex Addr	247F	9343
x"00",	-- Hex Addr	2480	9344
x"00",	-- Hex Addr	2481	9345
x"00",	-- Hex Addr	2482	9346
x"00",	-- Hex Addr	2483	9347
x"00",	-- Hex Addr	2484	9348
x"00",	-- Hex Addr	2485	9349
x"00",	-- Hex Addr	2486	9350
x"00",	-- Hex Addr	2487	9351
x"00",	-- Hex Addr	2488	9352
x"00",	-- Hex Addr	2489	9353
x"00",	-- Hex Addr	248A	9354
x"00",	-- Hex Addr	248B	9355
x"00",	-- Hex Addr	248C	9356
x"00",	-- Hex Addr	248D	9357
x"00",	-- Hex Addr	248E	9358
x"00",	-- Hex Addr	248F	9359
x"00",	-- Hex Addr	2490	9360
x"00",	-- Hex Addr	2491	9361
x"00",	-- Hex Addr	2492	9362
x"00",	-- Hex Addr	2493	9363
x"00",	-- Hex Addr	2494	9364
x"00",	-- Hex Addr	2495	9365
x"00",	-- Hex Addr	2496	9366
x"00",	-- Hex Addr	2497	9367
x"00",	-- Hex Addr	2498	9368
x"00",	-- Hex Addr	2499	9369
x"00",	-- Hex Addr	249A	9370
x"00",	-- Hex Addr	249B	9371
x"00",	-- Hex Addr	249C	9372
x"00",	-- Hex Addr	249D	9373
x"00",	-- Hex Addr	249E	9374
x"00",	-- Hex Addr	249F	9375
x"00",	-- Hex Addr	24A0	9376
x"00",	-- Hex Addr	24A1	9377
x"00",	-- Hex Addr	24A2	9378
x"00",	-- Hex Addr	24A3	9379
x"00",	-- Hex Addr	24A4	9380
x"00",	-- Hex Addr	24A5	9381
x"00",	-- Hex Addr	24A6	9382
x"00",	-- Hex Addr	24A7	9383
x"00",	-- Hex Addr	24A8	9384
x"00",	-- Hex Addr	24A9	9385
x"00",	-- Hex Addr	24AA	9386
x"00",	-- Hex Addr	24AB	9387
x"00",	-- Hex Addr	24AC	9388
x"00",	-- Hex Addr	24AD	9389
x"00",	-- Hex Addr	24AE	9390
x"00",	-- Hex Addr	24AF	9391
x"00",	-- Hex Addr	24B0	9392
x"00",	-- Hex Addr	24B1	9393
x"00",	-- Hex Addr	24B2	9394
x"00",	-- Hex Addr	24B3	9395
x"00",	-- Hex Addr	24B4	9396
x"00",	-- Hex Addr	24B5	9397
x"00",	-- Hex Addr	24B6	9398
x"00",	-- Hex Addr	24B7	9399
x"00",	-- Hex Addr	24B8	9400
x"00",	-- Hex Addr	24B9	9401
x"00",	-- Hex Addr	24BA	9402
x"00",	-- Hex Addr	24BB	9403
x"00",	-- Hex Addr	24BC	9404
x"00",	-- Hex Addr	24BD	9405
x"00",	-- Hex Addr	24BE	9406
x"00",	-- Hex Addr	24BF	9407
x"00",	-- Hex Addr	24C0	9408
x"00",	-- Hex Addr	24C1	9409
x"00",	-- Hex Addr	24C2	9410
x"00",	-- Hex Addr	24C3	9411
x"00",	-- Hex Addr	24C4	9412
x"00",	-- Hex Addr	24C5	9413
x"00",	-- Hex Addr	24C6	9414
x"00",	-- Hex Addr	24C7	9415
x"00",	-- Hex Addr	24C8	9416
x"00",	-- Hex Addr	24C9	9417
x"00",	-- Hex Addr	24CA	9418
x"00",	-- Hex Addr	24CB	9419
x"00",	-- Hex Addr	24CC	9420
x"00",	-- Hex Addr	24CD	9421
x"00",	-- Hex Addr	24CE	9422
x"00",	-- Hex Addr	24CF	9423
x"00",	-- Hex Addr	24D0	9424
x"00",	-- Hex Addr	24D1	9425
x"00",	-- Hex Addr	24D2	9426
x"00",	-- Hex Addr	24D3	9427
x"00",	-- Hex Addr	24D4	9428
x"00",	-- Hex Addr	24D5	9429
x"00",	-- Hex Addr	24D6	9430
x"00",	-- Hex Addr	24D7	9431
x"00",	-- Hex Addr	24D8	9432
x"00",	-- Hex Addr	24D9	9433
x"00",	-- Hex Addr	24DA	9434
x"00",	-- Hex Addr	24DB	9435
x"00",	-- Hex Addr	24DC	9436
x"00",	-- Hex Addr	24DD	9437
x"00",	-- Hex Addr	24DE	9438
x"00",	-- Hex Addr	24DF	9439
x"00",	-- Hex Addr	24E0	9440
x"00",	-- Hex Addr	24E1	9441
x"00",	-- Hex Addr	24E2	9442
x"00",	-- Hex Addr	24E3	9443
x"00",	-- Hex Addr	24E4	9444
x"00",	-- Hex Addr	24E5	9445
x"00",	-- Hex Addr	24E6	9446
x"00",	-- Hex Addr	24E7	9447
x"00",	-- Hex Addr	24E8	9448
x"00",	-- Hex Addr	24E9	9449
x"00",	-- Hex Addr	24EA	9450
x"00",	-- Hex Addr	24EB	9451
x"00",	-- Hex Addr	24EC	9452
x"00",	-- Hex Addr	24ED	9453
x"00",	-- Hex Addr	24EE	9454
x"00",	-- Hex Addr	24EF	9455
x"00",	-- Hex Addr	24F0	9456
x"00",	-- Hex Addr	24F1	9457
x"00",	-- Hex Addr	24F2	9458
x"00",	-- Hex Addr	24F3	9459
x"00",	-- Hex Addr	24F4	9460
x"00",	-- Hex Addr	24F5	9461
x"00",	-- Hex Addr	24F6	9462
x"00",	-- Hex Addr	24F7	9463
x"00",	-- Hex Addr	24F8	9464
x"00",	-- Hex Addr	24F9	9465
x"00",	-- Hex Addr	24FA	9466
x"00",	-- Hex Addr	24FB	9467
x"00",	-- Hex Addr	24FC	9468
x"00",	-- Hex Addr	24FD	9469
x"00",	-- Hex Addr	24FE	9470
x"00",	-- Hex Addr	24FF	9471
x"00",	-- Hex Addr	2500	9472
x"00",	-- Hex Addr	2501	9473
x"00",	-- Hex Addr	2502	9474
x"00",	-- Hex Addr	2503	9475
x"00",	-- Hex Addr	2504	9476
x"00",	-- Hex Addr	2505	9477
x"00",	-- Hex Addr	2506	9478
x"00",	-- Hex Addr	2507	9479
x"00",	-- Hex Addr	2508	9480
x"00",	-- Hex Addr	2509	9481
x"00",	-- Hex Addr	250A	9482
x"00",	-- Hex Addr	250B	9483
x"00",	-- Hex Addr	250C	9484
x"00",	-- Hex Addr	250D	9485
x"00",	-- Hex Addr	250E	9486
x"00",	-- Hex Addr	250F	9487
x"00",	-- Hex Addr	2510	9488
x"00",	-- Hex Addr	2511	9489
x"00",	-- Hex Addr	2512	9490
x"00",	-- Hex Addr	2513	9491
x"00",	-- Hex Addr	2514	9492
x"00",	-- Hex Addr	2515	9493
x"00",	-- Hex Addr	2516	9494
x"00",	-- Hex Addr	2517	9495
x"00",	-- Hex Addr	2518	9496
x"00",	-- Hex Addr	2519	9497
x"00",	-- Hex Addr	251A	9498
x"00",	-- Hex Addr	251B	9499
x"00",	-- Hex Addr	251C	9500
x"00",	-- Hex Addr	251D	9501
x"00",	-- Hex Addr	251E	9502
x"00",	-- Hex Addr	251F	9503
x"00",	-- Hex Addr	2520	9504
x"00",	-- Hex Addr	2521	9505
x"00",	-- Hex Addr	2522	9506
x"00",	-- Hex Addr	2523	9507
x"00",	-- Hex Addr	2524	9508
x"00",	-- Hex Addr	2525	9509
x"00",	-- Hex Addr	2526	9510
x"00",	-- Hex Addr	2527	9511
x"00",	-- Hex Addr	2528	9512
x"00",	-- Hex Addr	2529	9513
x"00",	-- Hex Addr	252A	9514
x"00",	-- Hex Addr	252B	9515
x"00",	-- Hex Addr	252C	9516
x"00",	-- Hex Addr	252D	9517
x"00",	-- Hex Addr	252E	9518
x"00",	-- Hex Addr	252F	9519
x"00",	-- Hex Addr	2530	9520
x"00",	-- Hex Addr	2531	9521
x"00",	-- Hex Addr	2532	9522
x"00",	-- Hex Addr	2533	9523
x"00",	-- Hex Addr	2534	9524
x"00",	-- Hex Addr	2535	9525
x"00",	-- Hex Addr	2536	9526
x"00",	-- Hex Addr	2537	9527
x"00",	-- Hex Addr	2538	9528
x"00",	-- Hex Addr	2539	9529
x"00",	-- Hex Addr	253A	9530
x"00",	-- Hex Addr	253B	9531
x"00",	-- Hex Addr	253C	9532
x"00",	-- Hex Addr	253D	9533
x"00",	-- Hex Addr	253E	9534
x"00",	-- Hex Addr	253F	9535
x"00",	-- Hex Addr	2540	9536
x"00",	-- Hex Addr	2541	9537
x"00",	-- Hex Addr	2542	9538
x"00",	-- Hex Addr	2543	9539
x"00",	-- Hex Addr	2544	9540
x"00",	-- Hex Addr	2545	9541
x"00",	-- Hex Addr	2546	9542
x"00",	-- Hex Addr	2547	9543
x"00",	-- Hex Addr	2548	9544
x"00",	-- Hex Addr	2549	9545
x"00",	-- Hex Addr	254A	9546
x"00",	-- Hex Addr	254B	9547
x"00",	-- Hex Addr	254C	9548
x"00",	-- Hex Addr	254D	9549
x"00",	-- Hex Addr	254E	9550
x"00",	-- Hex Addr	254F	9551
x"00",	-- Hex Addr	2550	9552
x"00",	-- Hex Addr	2551	9553
x"00",	-- Hex Addr	2552	9554
x"00",	-- Hex Addr	2553	9555
x"00",	-- Hex Addr	2554	9556
x"00",	-- Hex Addr	2555	9557
x"00",	-- Hex Addr	2556	9558
x"00",	-- Hex Addr	2557	9559
x"00",	-- Hex Addr	2558	9560
x"00",	-- Hex Addr	2559	9561
x"00",	-- Hex Addr	255A	9562
x"00",	-- Hex Addr	255B	9563
x"00",	-- Hex Addr	255C	9564
x"00",	-- Hex Addr	255D	9565
x"00",	-- Hex Addr	255E	9566
x"00",	-- Hex Addr	255F	9567
x"00",	-- Hex Addr	2560	9568
x"00",	-- Hex Addr	2561	9569
x"00",	-- Hex Addr	2562	9570
x"00",	-- Hex Addr	2563	9571
x"00",	-- Hex Addr	2564	9572
x"00",	-- Hex Addr	2565	9573
x"00",	-- Hex Addr	2566	9574
x"00",	-- Hex Addr	2567	9575
x"00",	-- Hex Addr	2568	9576
x"00",	-- Hex Addr	2569	9577
x"00",	-- Hex Addr	256A	9578
x"00",	-- Hex Addr	256B	9579
x"00",	-- Hex Addr	256C	9580
x"00",	-- Hex Addr	256D	9581
x"00",	-- Hex Addr	256E	9582
x"00",	-- Hex Addr	256F	9583
x"00",	-- Hex Addr	2570	9584
x"00",	-- Hex Addr	2571	9585
x"00",	-- Hex Addr	2572	9586
x"00",	-- Hex Addr	2573	9587
x"00",	-- Hex Addr	2574	9588
x"00",	-- Hex Addr	2575	9589
x"00",	-- Hex Addr	2576	9590
x"00",	-- Hex Addr	2577	9591
x"00",	-- Hex Addr	2578	9592
x"00",	-- Hex Addr	2579	9593
x"00",	-- Hex Addr	257A	9594
x"00",	-- Hex Addr	257B	9595
x"00",	-- Hex Addr	257C	9596
x"00",	-- Hex Addr	257D	9597
x"00",	-- Hex Addr	257E	9598
x"00",	-- Hex Addr	257F	9599
x"00",	-- Hex Addr	2580	9600
x"00",	-- Hex Addr	2581	9601
x"00",	-- Hex Addr	2582	9602
x"00",	-- Hex Addr	2583	9603
x"00",	-- Hex Addr	2584	9604
x"00",	-- Hex Addr	2585	9605
x"00",	-- Hex Addr	2586	9606
x"00",	-- Hex Addr	2587	9607
x"00",	-- Hex Addr	2588	9608
x"00",	-- Hex Addr	2589	9609
x"00",	-- Hex Addr	258A	9610
x"00",	-- Hex Addr	258B	9611
x"00",	-- Hex Addr	258C	9612
x"00",	-- Hex Addr	258D	9613
x"00",	-- Hex Addr	258E	9614
x"00",	-- Hex Addr	258F	9615
x"00",	-- Hex Addr	2590	9616
x"00",	-- Hex Addr	2591	9617
x"00",	-- Hex Addr	2592	9618
x"00",	-- Hex Addr	2593	9619
x"00",	-- Hex Addr	2594	9620
x"00",	-- Hex Addr	2595	9621
x"00",	-- Hex Addr	2596	9622
x"00",	-- Hex Addr	2597	9623
x"00",	-- Hex Addr	2598	9624
x"00",	-- Hex Addr	2599	9625
x"00",	-- Hex Addr	259A	9626
x"00",	-- Hex Addr	259B	9627
x"00",	-- Hex Addr	259C	9628
x"00",	-- Hex Addr	259D	9629
x"00",	-- Hex Addr	259E	9630
x"00",	-- Hex Addr	259F	9631
x"00",	-- Hex Addr	25A0	9632
x"00",	-- Hex Addr	25A1	9633
x"00",	-- Hex Addr	25A2	9634
x"00",	-- Hex Addr	25A3	9635
x"00",	-- Hex Addr	25A4	9636
x"00",	-- Hex Addr	25A5	9637
x"00",	-- Hex Addr	25A6	9638
x"00",	-- Hex Addr	25A7	9639
x"00",	-- Hex Addr	25A8	9640
x"00",	-- Hex Addr	25A9	9641
x"00",	-- Hex Addr	25AA	9642
x"00",	-- Hex Addr	25AB	9643
x"00",	-- Hex Addr	25AC	9644
x"00",	-- Hex Addr	25AD	9645
x"00",	-- Hex Addr	25AE	9646
x"00",	-- Hex Addr	25AF	9647
x"00",	-- Hex Addr	25B0	9648
x"00",	-- Hex Addr	25B1	9649
x"00",	-- Hex Addr	25B2	9650
x"00",	-- Hex Addr	25B3	9651
x"00",	-- Hex Addr	25B4	9652
x"00",	-- Hex Addr	25B5	9653
x"00",	-- Hex Addr	25B6	9654
x"00",	-- Hex Addr	25B7	9655
x"00",	-- Hex Addr	25B8	9656
x"00",	-- Hex Addr	25B9	9657
x"00",	-- Hex Addr	25BA	9658
x"00",	-- Hex Addr	25BB	9659
x"00",	-- Hex Addr	25BC	9660
x"00",	-- Hex Addr	25BD	9661
x"00",	-- Hex Addr	25BE	9662
x"00",	-- Hex Addr	25BF	9663
x"00",	-- Hex Addr	25C0	9664
x"00",	-- Hex Addr	25C1	9665
x"00",	-- Hex Addr	25C2	9666
x"00",	-- Hex Addr	25C3	9667
x"00",	-- Hex Addr	25C4	9668
x"00",	-- Hex Addr	25C5	9669
x"00",	-- Hex Addr	25C6	9670
x"00",	-- Hex Addr	25C7	9671
x"00",	-- Hex Addr	25C8	9672
x"00",	-- Hex Addr	25C9	9673
x"00",	-- Hex Addr	25CA	9674
x"00",	-- Hex Addr	25CB	9675
x"00",	-- Hex Addr	25CC	9676
x"00",	-- Hex Addr	25CD	9677
x"00",	-- Hex Addr	25CE	9678
x"00",	-- Hex Addr	25CF	9679
x"00",	-- Hex Addr	25D0	9680
x"00",	-- Hex Addr	25D1	9681
x"00",	-- Hex Addr	25D2	9682
x"00",	-- Hex Addr	25D3	9683
x"00",	-- Hex Addr	25D4	9684
x"00",	-- Hex Addr	25D5	9685
x"00",	-- Hex Addr	25D6	9686
x"00",	-- Hex Addr	25D7	9687
x"00",	-- Hex Addr	25D8	9688
x"00",	-- Hex Addr	25D9	9689
x"00",	-- Hex Addr	25DA	9690
x"00",	-- Hex Addr	25DB	9691
x"00",	-- Hex Addr	25DC	9692
x"00",	-- Hex Addr	25DD	9693
x"00",	-- Hex Addr	25DE	9694
x"00",	-- Hex Addr	25DF	9695
x"00",	-- Hex Addr	25E0	9696
x"00",	-- Hex Addr	25E1	9697
x"00",	-- Hex Addr	25E2	9698
x"00",	-- Hex Addr	25E3	9699
x"00",	-- Hex Addr	25E4	9700
x"00",	-- Hex Addr	25E5	9701
x"00",	-- Hex Addr	25E6	9702
x"00",	-- Hex Addr	25E7	9703
x"00",	-- Hex Addr	25E8	9704
x"00",	-- Hex Addr	25E9	9705
x"00",	-- Hex Addr	25EA	9706
x"00",	-- Hex Addr	25EB	9707
x"00",	-- Hex Addr	25EC	9708
x"00",	-- Hex Addr	25ED	9709
x"00",	-- Hex Addr	25EE	9710
x"00",	-- Hex Addr	25EF	9711
x"00",	-- Hex Addr	25F0	9712
x"00",	-- Hex Addr	25F1	9713
x"00",	-- Hex Addr	25F2	9714
x"00",	-- Hex Addr	25F3	9715
x"00",	-- Hex Addr	25F4	9716
x"00",	-- Hex Addr	25F5	9717
x"00",	-- Hex Addr	25F6	9718
x"00",	-- Hex Addr	25F7	9719
x"00",	-- Hex Addr	25F8	9720
x"00",	-- Hex Addr	25F9	9721
x"00",	-- Hex Addr	25FA	9722
x"00",	-- Hex Addr	25FB	9723
x"00",	-- Hex Addr	25FC	9724
x"00",	-- Hex Addr	25FD	9725
x"00",	-- Hex Addr	25FE	9726
x"00",	-- Hex Addr	25FF	9727
x"00",	-- Hex Addr	2600	9728
x"00",	-- Hex Addr	2601	9729
x"00",	-- Hex Addr	2602	9730
x"00",	-- Hex Addr	2603	9731
x"00",	-- Hex Addr	2604	9732
x"00",	-- Hex Addr	2605	9733
x"00",	-- Hex Addr	2606	9734
x"00",	-- Hex Addr	2607	9735
x"00",	-- Hex Addr	2608	9736
x"00",	-- Hex Addr	2609	9737
x"00",	-- Hex Addr	260A	9738
x"00",	-- Hex Addr	260B	9739
x"00",	-- Hex Addr	260C	9740
x"00",	-- Hex Addr	260D	9741
x"00",	-- Hex Addr	260E	9742
x"00",	-- Hex Addr	260F	9743
x"00",	-- Hex Addr	2610	9744
x"00",	-- Hex Addr	2611	9745
x"00",	-- Hex Addr	2612	9746
x"00",	-- Hex Addr	2613	9747
x"00",	-- Hex Addr	2614	9748
x"00",	-- Hex Addr	2615	9749
x"00",	-- Hex Addr	2616	9750
x"00",	-- Hex Addr	2617	9751
x"00",	-- Hex Addr	2618	9752
x"00",	-- Hex Addr	2619	9753
x"00",	-- Hex Addr	261A	9754
x"00",	-- Hex Addr	261B	9755
x"00",	-- Hex Addr	261C	9756
x"00",	-- Hex Addr	261D	9757
x"00",	-- Hex Addr	261E	9758
x"00",	-- Hex Addr	261F	9759
x"00",	-- Hex Addr	2620	9760
x"00",	-- Hex Addr	2621	9761
x"00",	-- Hex Addr	2622	9762
x"00",	-- Hex Addr	2623	9763
x"00",	-- Hex Addr	2624	9764
x"00",	-- Hex Addr	2625	9765
x"00",	-- Hex Addr	2626	9766
x"00",	-- Hex Addr	2627	9767
x"00",	-- Hex Addr	2628	9768
x"00",	-- Hex Addr	2629	9769
x"00",	-- Hex Addr	262A	9770
x"00",	-- Hex Addr	262B	9771
x"00",	-- Hex Addr	262C	9772
x"00",	-- Hex Addr	262D	9773
x"00",	-- Hex Addr	262E	9774
x"00",	-- Hex Addr	262F	9775
x"00",	-- Hex Addr	2630	9776
x"00",	-- Hex Addr	2631	9777
x"00",	-- Hex Addr	2632	9778
x"00",	-- Hex Addr	2633	9779
x"00",	-- Hex Addr	2634	9780
x"00",	-- Hex Addr	2635	9781
x"00",	-- Hex Addr	2636	9782
x"00",	-- Hex Addr	2637	9783
x"00",	-- Hex Addr	2638	9784
x"00",	-- Hex Addr	2639	9785
x"00",	-- Hex Addr	263A	9786
x"00",	-- Hex Addr	263B	9787
x"00",	-- Hex Addr	263C	9788
x"00",	-- Hex Addr	263D	9789
x"00",	-- Hex Addr	263E	9790
x"00",	-- Hex Addr	263F	9791
x"00",	-- Hex Addr	2640	9792
x"00",	-- Hex Addr	2641	9793
x"00",	-- Hex Addr	2642	9794
x"00",	-- Hex Addr	2643	9795
x"00",	-- Hex Addr	2644	9796
x"00",	-- Hex Addr	2645	9797
x"00",	-- Hex Addr	2646	9798
x"00",	-- Hex Addr	2647	9799
x"00",	-- Hex Addr	2648	9800
x"00",	-- Hex Addr	2649	9801
x"00",	-- Hex Addr	264A	9802
x"00",	-- Hex Addr	264B	9803
x"00",	-- Hex Addr	264C	9804
x"00",	-- Hex Addr	264D	9805
x"00",	-- Hex Addr	264E	9806
x"00",	-- Hex Addr	264F	9807
x"00",	-- Hex Addr	2650	9808
x"00",	-- Hex Addr	2651	9809
x"00",	-- Hex Addr	2652	9810
x"00",	-- Hex Addr	2653	9811
x"00",	-- Hex Addr	2654	9812
x"00",	-- Hex Addr	2655	9813
x"00",	-- Hex Addr	2656	9814
x"00",	-- Hex Addr	2657	9815
x"00",	-- Hex Addr	2658	9816
x"00",	-- Hex Addr	2659	9817
x"00",	-- Hex Addr	265A	9818
x"00",	-- Hex Addr	265B	9819
x"00",	-- Hex Addr	265C	9820
x"00",	-- Hex Addr	265D	9821
x"00",	-- Hex Addr	265E	9822
x"00",	-- Hex Addr	265F	9823
x"00",	-- Hex Addr	2660	9824
x"00",	-- Hex Addr	2661	9825
x"00",	-- Hex Addr	2662	9826
x"00",	-- Hex Addr	2663	9827
x"00",	-- Hex Addr	2664	9828
x"00",	-- Hex Addr	2665	9829
x"00",	-- Hex Addr	2666	9830
x"00",	-- Hex Addr	2667	9831
x"00",	-- Hex Addr	2668	9832
x"00",	-- Hex Addr	2669	9833
x"00",	-- Hex Addr	266A	9834
x"00",	-- Hex Addr	266B	9835
x"00",	-- Hex Addr	266C	9836
x"00",	-- Hex Addr	266D	9837
x"00",	-- Hex Addr	266E	9838
x"00",	-- Hex Addr	266F	9839
x"00",	-- Hex Addr	2670	9840
x"00",	-- Hex Addr	2671	9841
x"00",	-- Hex Addr	2672	9842
x"00",	-- Hex Addr	2673	9843
x"00",	-- Hex Addr	2674	9844
x"00",	-- Hex Addr	2675	9845
x"00",	-- Hex Addr	2676	9846
x"00",	-- Hex Addr	2677	9847
x"00",	-- Hex Addr	2678	9848
x"00",	-- Hex Addr	2679	9849
x"00",	-- Hex Addr	267A	9850
x"00",	-- Hex Addr	267B	9851
x"00",	-- Hex Addr	267C	9852
x"00",	-- Hex Addr	267D	9853
x"00",	-- Hex Addr	267E	9854
x"00",	-- Hex Addr	267F	9855
x"00",	-- Hex Addr	2680	9856
x"00",	-- Hex Addr	2681	9857
x"00",	-- Hex Addr	2682	9858
x"00",	-- Hex Addr	2683	9859
x"00",	-- Hex Addr	2684	9860
x"00",	-- Hex Addr	2685	9861
x"00",	-- Hex Addr	2686	9862
x"00",	-- Hex Addr	2687	9863
x"00",	-- Hex Addr	2688	9864
x"00",	-- Hex Addr	2689	9865
x"00",	-- Hex Addr	268A	9866
x"00",	-- Hex Addr	268B	9867
x"00",	-- Hex Addr	268C	9868
x"00",	-- Hex Addr	268D	9869
x"00",	-- Hex Addr	268E	9870
x"00",	-- Hex Addr	268F	9871
x"00",	-- Hex Addr	2690	9872
x"00",	-- Hex Addr	2691	9873
x"00",	-- Hex Addr	2692	9874
x"00",	-- Hex Addr	2693	9875
x"00",	-- Hex Addr	2694	9876
x"00",	-- Hex Addr	2695	9877
x"00",	-- Hex Addr	2696	9878
x"00",	-- Hex Addr	2697	9879
x"00",	-- Hex Addr	2698	9880
x"00",	-- Hex Addr	2699	9881
x"00",	-- Hex Addr	269A	9882
x"00",	-- Hex Addr	269B	9883
x"00",	-- Hex Addr	269C	9884
x"00",	-- Hex Addr	269D	9885
x"00",	-- Hex Addr	269E	9886
x"00",	-- Hex Addr	269F	9887
x"00",	-- Hex Addr	26A0	9888
x"00",	-- Hex Addr	26A1	9889
x"00",	-- Hex Addr	26A2	9890
x"00",	-- Hex Addr	26A3	9891
x"00",	-- Hex Addr	26A4	9892
x"00",	-- Hex Addr	26A5	9893
x"00",	-- Hex Addr	26A6	9894
x"00",	-- Hex Addr	26A7	9895
x"00",	-- Hex Addr	26A8	9896
x"00",	-- Hex Addr	26A9	9897
x"00",	-- Hex Addr	26AA	9898
x"00",	-- Hex Addr	26AB	9899
x"00",	-- Hex Addr	26AC	9900
x"00",	-- Hex Addr	26AD	9901
x"00",	-- Hex Addr	26AE	9902
x"00",	-- Hex Addr	26AF	9903
x"00",	-- Hex Addr	26B0	9904
x"00",	-- Hex Addr	26B1	9905
x"00",	-- Hex Addr	26B2	9906
x"00",	-- Hex Addr	26B3	9907
x"00",	-- Hex Addr	26B4	9908
x"00",	-- Hex Addr	26B5	9909
x"00",	-- Hex Addr	26B6	9910
x"00",	-- Hex Addr	26B7	9911
x"00",	-- Hex Addr	26B8	9912
x"00",	-- Hex Addr	26B9	9913
x"00",	-- Hex Addr	26BA	9914
x"00",	-- Hex Addr	26BB	9915
x"00",	-- Hex Addr	26BC	9916
x"00",	-- Hex Addr	26BD	9917
x"00",	-- Hex Addr	26BE	9918
x"00",	-- Hex Addr	26BF	9919
x"00",	-- Hex Addr	26C0	9920
x"00",	-- Hex Addr	26C1	9921
x"00",	-- Hex Addr	26C2	9922
x"00",	-- Hex Addr	26C3	9923
x"00",	-- Hex Addr	26C4	9924
x"00",	-- Hex Addr	26C5	9925
x"00",	-- Hex Addr	26C6	9926
x"00",	-- Hex Addr	26C7	9927
x"00",	-- Hex Addr	26C8	9928
x"00",	-- Hex Addr	26C9	9929
x"00",	-- Hex Addr	26CA	9930
x"00",	-- Hex Addr	26CB	9931
x"00",	-- Hex Addr	26CC	9932
x"00",	-- Hex Addr	26CD	9933
x"00",	-- Hex Addr	26CE	9934
x"00",	-- Hex Addr	26CF	9935
x"00",	-- Hex Addr	26D0	9936
x"00",	-- Hex Addr	26D1	9937
x"00",	-- Hex Addr	26D2	9938
x"00",	-- Hex Addr	26D3	9939
x"00",	-- Hex Addr	26D4	9940
x"00",	-- Hex Addr	26D5	9941
x"00",	-- Hex Addr	26D6	9942
x"00",	-- Hex Addr	26D7	9943
x"00",	-- Hex Addr	26D8	9944
x"00",	-- Hex Addr	26D9	9945
x"00",	-- Hex Addr	26DA	9946
x"00",	-- Hex Addr	26DB	9947
x"00",	-- Hex Addr	26DC	9948
x"00",	-- Hex Addr	26DD	9949
x"00",	-- Hex Addr	26DE	9950
x"00",	-- Hex Addr	26DF	9951
x"00",	-- Hex Addr	26E0	9952
x"00",	-- Hex Addr	26E1	9953
x"00",	-- Hex Addr	26E2	9954
x"00",	-- Hex Addr	26E3	9955
x"00",	-- Hex Addr	26E4	9956
x"00",	-- Hex Addr	26E5	9957
x"00",	-- Hex Addr	26E6	9958
x"00",	-- Hex Addr	26E7	9959
x"00",	-- Hex Addr	26E8	9960
x"00",	-- Hex Addr	26E9	9961
x"00",	-- Hex Addr	26EA	9962
x"00",	-- Hex Addr	26EB	9963
x"00",	-- Hex Addr	26EC	9964
x"00",	-- Hex Addr	26ED	9965
x"00",	-- Hex Addr	26EE	9966
x"00",	-- Hex Addr	26EF	9967
x"00",	-- Hex Addr	26F0	9968
x"00",	-- Hex Addr	26F1	9969
x"00",	-- Hex Addr	26F2	9970
x"00",	-- Hex Addr	26F3	9971
x"00",	-- Hex Addr	26F4	9972
x"00",	-- Hex Addr	26F5	9973
x"00",	-- Hex Addr	26F6	9974
x"00",	-- Hex Addr	26F7	9975
x"00",	-- Hex Addr	26F8	9976
x"00",	-- Hex Addr	26F9	9977
x"00",	-- Hex Addr	26FA	9978
x"00",	-- Hex Addr	26FB	9979
x"00",	-- Hex Addr	26FC	9980
x"00",	-- Hex Addr	26FD	9981
x"00",	-- Hex Addr	26FE	9982
x"00",	-- Hex Addr	26FF	9983
x"00",	-- Hex Addr	2700	9984
x"00",	-- Hex Addr	2701	9985
x"00",	-- Hex Addr	2702	9986
x"00",	-- Hex Addr	2703	9987
x"00",	-- Hex Addr	2704	9988
x"00",	-- Hex Addr	2705	9989
x"00",	-- Hex Addr	2706	9990
x"00",	-- Hex Addr	2707	9991
x"00",	-- Hex Addr	2708	9992
x"00",	-- Hex Addr	2709	9993
x"00",	-- Hex Addr	270A	9994
x"00",	-- Hex Addr	270B	9995
x"00",	-- Hex Addr	270C	9996
x"00",	-- Hex Addr	270D	9997
x"00",	-- Hex Addr	270E	9998
x"00",	-- Hex Addr	270F	9999
x"00",	-- Hex Addr	2710	10000
x"00",	-- Hex Addr	2711	10001
x"00",	-- Hex Addr	2712	10002
x"00",	-- Hex Addr	2713	10003
x"00",	-- Hex Addr	2714	10004
x"00",	-- Hex Addr	2715	10005
x"00",	-- Hex Addr	2716	10006
x"00",	-- Hex Addr	2717	10007
x"00",	-- Hex Addr	2718	10008
x"00",	-- Hex Addr	2719	10009
x"00",	-- Hex Addr	271A	10010
x"00",	-- Hex Addr	271B	10011
x"00",	-- Hex Addr	271C	10012
x"00",	-- Hex Addr	271D	10013
x"00",	-- Hex Addr	271E	10014
x"00",	-- Hex Addr	271F	10015
x"00",	-- Hex Addr	2720	10016
x"00",	-- Hex Addr	2721	10017
x"00",	-- Hex Addr	2722	10018
x"00",	-- Hex Addr	2723	10019
x"00",	-- Hex Addr	2724	10020
x"00",	-- Hex Addr	2725	10021
x"00",	-- Hex Addr	2726	10022
x"00",	-- Hex Addr	2727	10023
x"00",	-- Hex Addr	2728	10024
x"00",	-- Hex Addr	2729	10025
x"00",	-- Hex Addr	272A	10026
x"00",	-- Hex Addr	272B	10027
x"00",	-- Hex Addr	272C	10028
x"00",	-- Hex Addr	272D	10029
x"00",	-- Hex Addr	272E	10030
x"00",	-- Hex Addr	272F	10031
x"00",	-- Hex Addr	2730	10032
x"00",	-- Hex Addr	2731	10033
x"00",	-- Hex Addr	2732	10034
x"00",	-- Hex Addr	2733	10035
x"00",	-- Hex Addr	2734	10036
x"00",	-- Hex Addr	2735	10037
x"00",	-- Hex Addr	2736	10038
x"00",	-- Hex Addr	2737	10039
x"00",	-- Hex Addr	2738	10040
x"00",	-- Hex Addr	2739	10041
x"00",	-- Hex Addr	273A	10042
x"00",	-- Hex Addr	273B	10043
x"00",	-- Hex Addr	273C	10044
x"00",	-- Hex Addr	273D	10045
x"00",	-- Hex Addr	273E	10046
x"00",	-- Hex Addr	273F	10047
x"00",	-- Hex Addr	2740	10048
x"00",	-- Hex Addr	2741	10049
x"00",	-- Hex Addr	2742	10050
x"00",	-- Hex Addr	2743	10051
x"00",	-- Hex Addr	2744	10052
x"00",	-- Hex Addr	2745	10053
x"00",	-- Hex Addr	2746	10054
x"00",	-- Hex Addr	2747	10055
x"00",	-- Hex Addr	2748	10056
x"00",	-- Hex Addr	2749	10057
x"00",	-- Hex Addr	274A	10058
x"00",	-- Hex Addr	274B	10059
x"00",	-- Hex Addr	274C	10060
x"00",	-- Hex Addr	274D	10061
x"00",	-- Hex Addr	274E	10062
x"00",	-- Hex Addr	274F	10063
x"00",	-- Hex Addr	2750	10064
x"00",	-- Hex Addr	2751	10065
x"00",	-- Hex Addr	2752	10066
x"00",	-- Hex Addr	2753	10067
x"00",	-- Hex Addr	2754	10068
x"00",	-- Hex Addr	2755	10069
x"00",	-- Hex Addr	2756	10070
x"00",	-- Hex Addr	2757	10071
x"00",	-- Hex Addr	2758	10072
x"00",	-- Hex Addr	2759	10073
x"00",	-- Hex Addr	275A	10074
x"00",	-- Hex Addr	275B	10075
x"00",	-- Hex Addr	275C	10076
x"00",	-- Hex Addr	275D	10077
x"00",	-- Hex Addr	275E	10078
x"00",	-- Hex Addr	275F	10079
x"00",	-- Hex Addr	2760	10080
x"00",	-- Hex Addr	2761	10081
x"00",	-- Hex Addr	2762	10082
x"00",	-- Hex Addr	2763	10083
x"00",	-- Hex Addr	2764	10084
x"00",	-- Hex Addr	2765	10085
x"00",	-- Hex Addr	2766	10086
x"00",	-- Hex Addr	2767	10087
x"00",	-- Hex Addr	2768	10088
x"00",	-- Hex Addr	2769	10089
x"00",	-- Hex Addr	276A	10090
x"00",	-- Hex Addr	276B	10091
x"00",	-- Hex Addr	276C	10092
x"00",	-- Hex Addr	276D	10093
x"00",	-- Hex Addr	276E	10094
x"00",	-- Hex Addr	276F	10095
x"00",	-- Hex Addr	2770	10096
x"00",	-- Hex Addr	2771	10097
x"00",	-- Hex Addr	2772	10098
x"00",	-- Hex Addr	2773	10099
x"00",	-- Hex Addr	2774	10100
x"00",	-- Hex Addr	2775	10101
x"00",	-- Hex Addr	2776	10102
x"00",	-- Hex Addr	2777	10103
x"00",	-- Hex Addr	2778	10104
x"00",	-- Hex Addr	2779	10105
x"00",	-- Hex Addr	277A	10106
x"00",	-- Hex Addr	277B	10107
x"00",	-- Hex Addr	277C	10108
x"00",	-- Hex Addr	277D	10109
x"00",	-- Hex Addr	277E	10110
x"00",	-- Hex Addr	277F	10111
x"00",	-- Hex Addr	2780	10112
x"00",	-- Hex Addr	2781	10113
x"00",	-- Hex Addr	2782	10114
x"00",	-- Hex Addr	2783	10115
x"00",	-- Hex Addr	2784	10116
x"00",	-- Hex Addr	2785	10117
x"00",	-- Hex Addr	2786	10118
x"00",	-- Hex Addr	2787	10119
x"00",	-- Hex Addr	2788	10120
x"00",	-- Hex Addr	2789	10121
x"00",	-- Hex Addr	278A	10122
x"00",	-- Hex Addr	278B	10123
x"00",	-- Hex Addr	278C	10124
x"00",	-- Hex Addr	278D	10125
x"00",	-- Hex Addr	278E	10126
x"00",	-- Hex Addr	278F	10127
x"00",	-- Hex Addr	2790	10128
x"00",	-- Hex Addr	2791	10129
x"00",	-- Hex Addr	2792	10130
x"00",	-- Hex Addr	2793	10131
x"00",	-- Hex Addr	2794	10132
x"00",	-- Hex Addr	2795	10133
x"00",	-- Hex Addr	2796	10134
x"00",	-- Hex Addr	2797	10135
x"00",	-- Hex Addr	2798	10136
x"00",	-- Hex Addr	2799	10137
x"00",	-- Hex Addr	279A	10138
x"00",	-- Hex Addr	279B	10139
x"00",	-- Hex Addr	279C	10140
x"00",	-- Hex Addr	279D	10141
x"00",	-- Hex Addr	279E	10142
x"00",	-- Hex Addr	279F	10143
x"00",	-- Hex Addr	27A0	10144
x"00",	-- Hex Addr	27A1	10145
x"00",	-- Hex Addr	27A2	10146
x"00",	-- Hex Addr	27A3	10147
x"00",	-- Hex Addr	27A4	10148
x"00",	-- Hex Addr	27A5	10149
x"00",	-- Hex Addr	27A6	10150
x"00",	-- Hex Addr	27A7	10151
x"00",	-- Hex Addr	27A8	10152
x"00",	-- Hex Addr	27A9	10153
x"00",	-- Hex Addr	27AA	10154
x"00",	-- Hex Addr	27AB	10155
x"00",	-- Hex Addr	27AC	10156
x"00",	-- Hex Addr	27AD	10157
x"00",	-- Hex Addr	27AE	10158
x"00",	-- Hex Addr	27AF	10159
x"00",	-- Hex Addr	27B0	10160
x"00",	-- Hex Addr	27B1	10161
x"00",	-- Hex Addr	27B2	10162
x"00",	-- Hex Addr	27B3	10163
x"00",	-- Hex Addr	27B4	10164
x"00",	-- Hex Addr	27B5	10165
x"00",	-- Hex Addr	27B6	10166
x"00",	-- Hex Addr	27B7	10167
x"00",	-- Hex Addr	27B8	10168
x"00",	-- Hex Addr	27B9	10169
x"00",	-- Hex Addr	27BA	10170
x"00",	-- Hex Addr	27BB	10171
x"00",	-- Hex Addr	27BC	10172
x"00",	-- Hex Addr	27BD	10173
x"00",	-- Hex Addr	27BE	10174
x"00",	-- Hex Addr	27BF	10175
x"00",	-- Hex Addr	27C0	10176
x"00",	-- Hex Addr	27C1	10177
x"00",	-- Hex Addr	27C2	10178
x"00",	-- Hex Addr	27C3	10179
x"00",	-- Hex Addr	27C4	10180
x"00",	-- Hex Addr	27C5	10181
x"00",	-- Hex Addr	27C6	10182
x"00",	-- Hex Addr	27C7	10183
x"00",	-- Hex Addr	27C8	10184
x"00",	-- Hex Addr	27C9	10185
x"00",	-- Hex Addr	27CA	10186
x"00",	-- Hex Addr	27CB	10187
x"00",	-- Hex Addr	27CC	10188
x"00",	-- Hex Addr	27CD	10189
x"00",	-- Hex Addr	27CE	10190
x"00",	-- Hex Addr	27CF	10191
x"00",	-- Hex Addr	27D0	10192
x"00",	-- Hex Addr	27D1	10193
x"00",	-- Hex Addr	27D2	10194
x"00",	-- Hex Addr	27D3	10195
x"00",	-- Hex Addr	27D4	10196
x"00",	-- Hex Addr	27D5	10197
x"00",	-- Hex Addr	27D6	10198
x"00",	-- Hex Addr	27D7	10199
x"00",	-- Hex Addr	27D8	10200
x"00",	-- Hex Addr	27D9	10201
x"00",	-- Hex Addr	27DA	10202
x"00",	-- Hex Addr	27DB	10203
x"00",	-- Hex Addr	27DC	10204
x"00",	-- Hex Addr	27DD	10205
x"00",	-- Hex Addr	27DE	10206
x"00",	-- Hex Addr	27DF	10207
x"00",	-- Hex Addr	27E0	10208
x"00",	-- Hex Addr	27E1	10209
x"00",	-- Hex Addr	27E2	10210
x"00",	-- Hex Addr	27E3	10211
x"00",	-- Hex Addr	27E4	10212
x"00",	-- Hex Addr	27E5	10213
x"00",	-- Hex Addr	27E6	10214
x"00",	-- Hex Addr	27E7	10215
x"00",	-- Hex Addr	27E8	10216
x"00",	-- Hex Addr	27E9	10217
x"00",	-- Hex Addr	27EA	10218
x"00",	-- Hex Addr	27EB	10219
x"00",	-- Hex Addr	27EC	10220
x"00",	-- Hex Addr	27ED	10221
x"00",	-- Hex Addr	27EE	10222
x"00",	-- Hex Addr	27EF	10223
x"00",	-- Hex Addr	27F0	10224
x"00",	-- Hex Addr	27F1	10225
x"00",	-- Hex Addr	27F2	10226
x"00",	-- Hex Addr	27F3	10227
x"00",	-- Hex Addr	27F4	10228
x"00",	-- Hex Addr	27F5	10229
x"00",	-- Hex Addr	27F6	10230
x"00",	-- Hex Addr	27F7	10231
x"00",	-- Hex Addr	27F8	10232
x"00",	-- Hex Addr	27F9	10233
x"00",	-- Hex Addr	27FA	10234
x"00",	-- Hex Addr	27FB	10235
x"00",	-- Hex Addr	27FC	10236
x"00",	-- Hex Addr	27FD	10237
x"00",	-- Hex Addr	27FE	10238
x"00",	-- Hex Addr	27FF	10239
x"00",	-- Hex Addr	2800	10240
x"00",	-- Hex Addr	2801	10241
x"00",	-- Hex Addr	2802	10242
x"00",	-- Hex Addr	2803	10243
x"00",	-- Hex Addr	2804	10244
x"00",	-- Hex Addr	2805	10245
x"00",	-- Hex Addr	2806	10246
x"00",	-- Hex Addr	2807	10247
x"00",	-- Hex Addr	2808	10248
x"00",	-- Hex Addr	2809	10249
x"00",	-- Hex Addr	280A	10250
x"00",	-- Hex Addr	280B	10251
x"00",	-- Hex Addr	280C	10252
x"00",	-- Hex Addr	280D	10253
x"00",	-- Hex Addr	280E	10254
x"00",	-- Hex Addr	280F	10255
x"00",	-- Hex Addr	2810	10256
x"00",	-- Hex Addr	2811	10257
x"00",	-- Hex Addr	2812	10258
x"00",	-- Hex Addr	2813	10259
x"00",	-- Hex Addr	2814	10260
x"00",	-- Hex Addr	2815	10261
x"00",	-- Hex Addr	2816	10262
x"00",	-- Hex Addr	2817	10263
x"00",	-- Hex Addr	2818	10264
x"00",	-- Hex Addr	2819	10265
x"00",	-- Hex Addr	281A	10266
x"00",	-- Hex Addr	281B	10267
x"00",	-- Hex Addr	281C	10268
x"00",	-- Hex Addr	281D	10269
x"00",	-- Hex Addr	281E	10270
x"00",	-- Hex Addr	281F	10271
x"00",	-- Hex Addr	2820	10272
x"00",	-- Hex Addr	2821	10273
x"00",	-- Hex Addr	2822	10274
x"00",	-- Hex Addr	2823	10275
x"00",	-- Hex Addr	2824	10276
x"00",	-- Hex Addr	2825	10277
x"00",	-- Hex Addr	2826	10278
x"00",	-- Hex Addr	2827	10279
x"00",	-- Hex Addr	2828	10280
x"00",	-- Hex Addr	2829	10281
x"00",	-- Hex Addr	282A	10282
x"00",	-- Hex Addr	282B	10283
x"00",	-- Hex Addr	282C	10284
x"00",	-- Hex Addr	282D	10285
x"00",	-- Hex Addr	282E	10286
x"00",	-- Hex Addr	282F	10287
x"00",	-- Hex Addr	2830	10288
x"00",	-- Hex Addr	2831	10289
x"00",	-- Hex Addr	2832	10290
x"00",	-- Hex Addr	2833	10291
x"00",	-- Hex Addr	2834	10292
x"00",	-- Hex Addr	2835	10293
x"00",	-- Hex Addr	2836	10294
x"00",	-- Hex Addr	2837	10295
x"00",	-- Hex Addr	2838	10296
x"00",	-- Hex Addr	2839	10297
x"00",	-- Hex Addr	283A	10298
x"00",	-- Hex Addr	283B	10299
x"00",	-- Hex Addr	283C	10300
x"00",	-- Hex Addr	283D	10301
x"00",	-- Hex Addr	283E	10302
x"00",	-- Hex Addr	283F	10303
x"00",	-- Hex Addr	2840	10304
x"00",	-- Hex Addr	2841	10305
x"00",	-- Hex Addr	2842	10306
x"00",	-- Hex Addr	2843	10307
x"00",	-- Hex Addr	2844	10308
x"00",	-- Hex Addr	2845	10309
x"00",	-- Hex Addr	2846	10310
x"00",	-- Hex Addr	2847	10311
x"00",	-- Hex Addr	2848	10312
x"00",	-- Hex Addr	2849	10313
x"00",	-- Hex Addr	284A	10314
x"00",	-- Hex Addr	284B	10315
x"00",	-- Hex Addr	284C	10316
x"00",	-- Hex Addr	284D	10317
x"00",	-- Hex Addr	284E	10318
x"00",	-- Hex Addr	284F	10319
x"00",	-- Hex Addr	2850	10320
x"00",	-- Hex Addr	2851	10321
x"00",	-- Hex Addr	2852	10322
x"00",	-- Hex Addr	2853	10323
x"00",	-- Hex Addr	2854	10324
x"00",	-- Hex Addr	2855	10325
x"00",	-- Hex Addr	2856	10326
x"00",	-- Hex Addr	2857	10327
x"00",	-- Hex Addr	2858	10328
x"00",	-- Hex Addr	2859	10329
x"00",	-- Hex Addr	285A	10330
x"00",	-- Hex Addr	285B	10331
x"00",	-- Hex Addr	285C	10332
x"00",	-- Hex Addr	285D	10333
x"00",	-- Hex Addr	285E	10334
x"00",	-- Hex Addr	285F	10335
x"00",	-- Hex Addr	2860	10336
x"00",	-- Hex Addr	2861	10337
x"00",	-- Hex Addr	2862	10338
x"00",	-- Hex Addr	2863	10339
x"00",	-- Hex Addr	2864	10340
x"00",	-- Hex Addr	2865	10341
x"00",	-- Hex Addr	2866	10342
x"00",	-- Hex Addr	2867	10343
x"00",	-- Hex Addr	2868	10344
x"00",	-- Hex Addr	2869	10345
x"00",	-- Hex Addr	286A	10346
x"00",	-- Hex Addr	286B	10347
x"00",	-- Hex Addr	286C	10348
x"00",	-- Hex Addr	286D	10349
x"00",	-- Hex Addr	286E	10350
x"00",	-- Hex Addr	286F	10351
x"00",	-- Hex Addr	2870	10352
x"00",	-- Hex Addr	2871	10353
x"00",	-- Hex Addr	2872	10354
x"00",	-- Hex Addr	2873	10355
x"00",	-- Hex Addr	2874	10356
x"00",	-- Hex Addr	2875	10357
x"00",	-- Hex Addr	2876	10358
x"00",	-- Hex Addr	2877	10359
x"00",	-- Hex Addr	2878	10360
x"00",	-- Hex Addr	2879	10361
x"00",	-- Hex Addr	287A	10362
x"00",	-- Hex Addr	287B	10363
x"00",	-- Hex Addr	287C	10364
x"00",	-- Hex Addr	287D	10365
x"00",	-- Hex Addr	287E	10366
x"00",	-- Hex Addr	287F	10367
x"00",	-- Hex Addr	2880	10368
x"00",	-- Hex Addr	2881	10369
x"00",	-- Hex Addr	2882	10370
x"00",	-- Hex Addr	2883	10371
x"00",	-- Hex Addr	2884	10372
x"00",	-- Hex Addr	2885	10373
x"00",	-- Hex Addr	2886	10374
x"00",	-- Hex Addr	2887	10375
x"00",	-- Hex Addr	2888	10376
x"00",	-- Hex Addr	2889	10377
x"00",	-- Hex Addr	288A	10378
x"00",	-- Hex Addr	288B	10379
x"00",	-- Hex Addr	288C	10380
x"00",	-- Hex Addr	288D	10381
x"00",	-- Hex Addr	288E	10382
x"00",	-- Hex Addr	288F	10383
x"00",	-- Hex Addr	2890	10384
x"00",	-- Hex Addr	2891	10385
x"00",	-- Hex Addr	2892	10386
x"00",	-- Hex Addr	2893	10387
x"00",	-- Hex Addr	2894	10388
x"00",	-- Hex Addr	2895	10389
x"00",	-- Hex Addr	2896	10390
x"00",	-- Hex Addr	2897	10391
x"00",	-- Hex Addr	2898	10392
x"00",	-- Hex Addr	2899	10393
x"00",	-- Hex Addr	289A	10394
x"00",	-- Hex Addr	289B	10395
x"00",	-- Hex Addr	289C	10396
x"00",	-- Hex Addr	289D	10397
x"00",	-- Hex Addr	289E	10398
x"00",	-- Hex Addr	289F	10399
x"00",	-- Hex Addr	28A0	10400
x"00",	-- Hex Addr	28A1	10401
x"00",	-- Hex Addr	28A2	10402
x"00",	-- Hex Addr	28A3	10403
x"00",	-- Hex Addr	28A4	10404
x"00",	-- Hex Addr	28A5	10405
x"00",	-- Hex Addr	28A6	10406
x"00",	-- Hex Addr	28A7	10407
x"00",	-- Hex Addr	28A8	10408
x"00",	-- Hex Addr	28A9	10409
x"00",	-- Hex Addr	28AA	10410
x"00",	-- Hex Addr	28AB	10411
x"00",	-- Hex Addr	28AC	10412
x"00",	-- Hex Addr	28AD	10413
x"00",	-- Hex Addr	28AE	10414
x"00",	-- Hex Addr	28AF	10415
x"00",	-- Hex Addr	28B0	10416
x"00",	-- Hex Addr	28B1	10417
x"00",	-- Hex Addr	28B2	10418
x"00",	-- Hex Addr	28B3	10419
x"00",	-- Hex Addr	28B4	10420
x"00",	-- Hex Addr	28B5	10421
x"00",	-- Hex Addr	28B6	10422
x"00",	-- Hex Addr	28B7	10423
x"00",	-- Hex Addr	28B8	10424
x"00",	-- Hex Addr	28B9	10425
x"00",	-- Hex Addr	28BA	10426
x"00",	-- Hex Addr	28BB	10427
x"00",	-- Hex Addr	28BC	10428
x"00",	-- Hex Addr	28BD	10429
x"00",	-- Hex Addr	28BE	10430
x"00",	-- Hex Addr	28BF	10431
x"00",	-- Hex Addr	28C0	10432
x"00",	-- Hex Addr	28C1	10433
x"00",	-- Hex Addr	28C2	10434
x"00",	-- Hex Addr	28C3	10435
x"00",	-- Hex Addr	28C4	10436
x"00",	-- Hex Addr	28C5	10437
x"00",	-- Hex Addr	28C6	10438
x"00",	-- Hex Addr	28C7	10439
x"00",	-- Hex Addr	28C8	10440
x"00",	-- Hex Addr	28C9	10441
x"00",	-- Hex Addr	28CA	10442
x"00",	-- Hex Addr	28CB	10443
x"00",	-- Hex Addr	28CC	10444
x"00",	-- Hex Addr	28CD	10445
x"00",	-- Hex Addr	28CE	10446
x"00",	-- Hex Addr	28CF	10447
x"00",	-- Hex Addr	28D0	10448
x"00",	-- Hex Addr	28D1	10449
x"00",	-- Hex Addr	28D2	10450
x"00",	-- Hex Addr	28D3	10451
x"00",	-- Hex Addr	28D4	10452
x"00",	-- Hex Addr	28D5	10453
x"00",	-- Hex Addr	28D6	10454
x"00",	-- Hex Addr	28D7	10455
x"00",	-- Hex Addr	28D8	10456
x"00",	-- Hex Addr	28D9	10457
x"00",	-- Hex Addr	28DA	10458
x"00",	-- Hex Addr	28DB	10459
x"00",	-- Hex Addr	28DC	10460
x"00",	-- Hex Addr	28DD	10461
x"00",	-- Hex Addr	28DE	10462
x"00",	-- Hex Addr	28DF	10463
x"00",	-- Hex Addr	28E0	10464
x"00",	-- Hex Addr	28E1	10465
x"00",	-- Hex Addr	28E2	10466
x"00",	-- Hex Addr	28E3	10467
x"00",	-- Hex Addr	28E4	10468
x"00",	-- Hex Addr	28E5	10469
x"00",	-- Hex Addr	28E6	10470
x"00",	-- Hex Addr	28E7	10471
x"00",	-- Hex Addr	28E8	10472
x"00",	-- Hex Addr	28E9	10473
x"00",	-- Hex Addr	28EA	10474
x"00",	-- Hex Addr	28EB	10475
x"00",	-- Hex Addr	28EC	10476
x"00",	-- Hex Addr	28ED	10477
x"00",	-- Hex Addr	28EE	10478
x"00",	-- Hex Addr	28EF	10479
x"00",	-- Hex Addr	28F0	10480
x"00",	-- Hex Addr	28F1	10481
x"00",	-- Hex Addr	28F2	10482
x"00",	-- Hex Addr	28F3	10483
x"00",	-- Hex Addr	28F4	10484
x"00",	-- Hex Addr	28F5	10485
x"00",	-- Hex Addr	28F6	10486
x"00",	-- Hex Addr	28F7	10487
x"00",	-- Hex Addr	28F8	10488
x"00",	-- Hex Addr	28F9	10489
x"00",	-- Hex Addr	28FA	10490
x"00",	-- Hex Addr	28FB	10491
x"00",	-- Hex Addr	28FC	10492
x"00",	-- Hex Addr	28FD	10493
x"00",	-- Hex Addr	28FE	10494
x"00",	-- Hex Addr	28FF	10495
x"00",	-- Hex Addr	2900	10496
x"00",	-- Hex Addr	2901	10497
x"00",	-- Hex Addr	2902	10498
x"00",	-- Hex Addr	2903	10499
x"00",	-- Hex Addr	2904	10500
x"00",	-- Hex Addr	2905	10501
x"00",	-- Hex Addr	2906	10502
x"00",	-- Hex Addr	2907	10503
x"00",	-- Hex Addr	2908	10504
x"00",	-- Hex Addr	2909	10505
x"00",	-- Hex Addr	290A	10506
x"00",	-- Hex Addr	290B	10507
x"00",	-- Hex Addr	290C	10508
x"00",	-- Hex Addr	290D	10509
x"00",	-- Hex Addr	290E	10510
x"00",	-- Hex Addr	290F	10511
x"00",	-- Hex Addr	2910	10512
x"00",	-- Hex Addr	2911	10513
x"00",	-- Hex Addr	2912	10514
x"00",	-- Hex Addr	2913	10515
x"00",	-- Hex Addr	2914	10516
x"00",	-- Hex Addr	2915	10517
x"00",	-- Hex Addr	2916	10518
x"00",	-- Hex Addr	2917	10519
x"00",	-- Hex Addr	2918	10520
x"00",	-- Hex Addr	2919	10521
x"00",	-- Hex Addr	291A	10522
x"00",	-- Hex Addr	291B	10523
x"00",	-- Hex Addr	291C	10524
x"00",	-- Hex Addr	291D	10525
x"00",	-- Hex Addr	291E	10526
x"00",	-- Hex Addr	291F	10527
x"00",	-- Hex Addr	2920	10528
x"00",	-- Hex Addr	2921	10529
x"00",	-- Hex Addr	2922	10530
x"00",	-- Hex Addr	2923	10531
x"00",	-- Hex Addr	2924	10532
x"00",	-- Hex Addr	2925	10533
x"00",	-- Hex Addr	2926	10534
x"00",	-- Hex Addr	2927	10535
x"00",	-- Hex Addr	2928	10536
x"00",	-- Hex Addr	2929	10537
x"00",	-- Hex Addr	292A	10538
x"00",	-- Hex Addr	292B	10539
x"00",	-- Hex Addr	292C	10540
x"00",	-- Hex Addr	292D	10541
x"00",	-- Hex Addr	292E	10542
x"00",	-- Hex Addr	292F	10543
x"00",	-- Hex Addr	2930	10544
x"00",	-- Hex Addr	2931	10545
x"00",	-- Hex Addr	2932	10546
x"00",	-- Hex Addr	2933	10547
x"00",	-- Hex Addr	2934	10548
x"00",	-- Hex Addr	2935	10549
x"00",	-- Hex Addr	2936	10550
x"00",	-- Hex Addr	2937	10551
x"00",	-- Hex Addr	2938	10552
x"00",	-- Hex Addr	2939	10553
x"00",	-- Hex Addr	293A	10554
x"00",	-- Hex Addr	293B	10555
x"00",	-- Hex Addr	293C	10556
x"00",	-- Hex Addr	293D	10557
x"00",	-- Hex Addr	293E	10558
x"00",	-- Hex Addr	293F	10559
x"00",	-- Hex Addr	2940	10560
x"00",	-- Hex Addr	2941	10561
x"00",	-- Hex Addr	2942	10562
x"00",	-- Hex Addr	2943	10563
x"00",	-- Hex Addr	2944	10564
x"00",	-- Hex Addr	2945	10565
x"00",	-- Hex Addr	2946	10566
x"00",	-- Hex Addr	2947	10567
x"00",	-- Hex Addr	2948	10568
x"00",	-- Hex Addr	2949	10569
x"00",	-- Hex Addr	294A	10570
x"00",	-- Hex Addr	294B	10571
x"00",	-- Hex Addr	294C	10572
x"00",	-- Hex Addr	294D	10573
x"00",	-- Hex Addr	294E	10574
x"00",	-- Hex Addr	294F	10575
x"00",	-- Hex Addr	2950	10576
x"00",	-- Hex Addr	2951	10577
x"00",	-- Hex Addr	2952	10578
x"00",	-- Hex Addr	2953	10579
x"00",	-- Hex Addr	2954	10580
x"00",	-- Hex Addr	2955	10581
x"00",	-- Hex Addr	2956	10582
x"00",	-- Hex Addr	2957	10583
x"00",	-- Hex Addr	2958	10584
x"00",	-- Hex Addr	2959	10585
x"00",	-- Hex Addr	295A	10586
x"00",	-- Hex Addr	295B	10587
x"00",	-- Hex Addr	295C	10588
x"00",	-- Hex Addr	295D	10589
x"00",	-- Hex Addr	295E	10590
x"00",	-- Hex Addr	295F	10591
x"00",	-- Hex Addr	2960	10592
x"00",	-- Hex Addr	2961	10593
x"00",	-- Hex Addr	2962	10594
x"00",	-- Hex Addr	2963	10595
x"00",	-- Hex Addr	2964	10596
x"00",	-- Hex Addr	2965	10597
x"00",	-- Hex Addr	2966	10598
x"00",	-- Hex Addr	2967	10599
x"00",	-- Hex Addr	2968	10600
x"00",	-- Hex Addr	2969	10601
x"00",	-- Hex Addr	296A	10602
x"00",	-- Hex Addr	296B	10603
x"00",	-- Hex Addr	296C	10604
x"00",	-- Hex Addr	296D	10605
x"00",	-- Hex Addr	296E	10606
x"00",	-- Hex Addr	296F	10607
x"00",	-- Hex Addr	2970	10608
x"00",	-- Hex Addr	2971	10609
x"00",	-- Hex Addr	2972	10610
x"00",	-- Hex Addr	2973	10611
x"00",	-- Hex Addr	2974	10612
x"00",	-- Hex Addr	2975	10613
x"00",	-- Hex Addr	2976	10614
x"00",	-- Hex Addr	2977	10615
x"00",	-- Hex Addr	2978	10616
x"00",	-- Hex Addr	2979	10617
x"00",	-- Hex Addr	297A	10618
x"00",	-- Hex Addr	297B	10619
x"00",	-- Hex Addr	297C	10620
x"00",	-- Hex Addr	297D	10621
x"00",	-- Hex Addr	297E	10622
x"00",	-- Hex Addr	297F	10623
x"00",	-- Hex Addr	2980	10624
x"00",	-- Hex Addr	2981	10625
x"00",	-- Hex Addr	2982	10626
x"00",	-- Hex Addr	2983	10627
x"00",	-- Hex Addr	2984	10628
x"00",	-- Hex Addr	2985	10629
x"00",	-- Hex Addr	2986	10630
x"00",	-- Hex Addr	2987	10631
x"00",	-- Hex Addr	2988	10632
x"00",	-- Hex Addr	2989	10633
x"00",	-- Hex Addr	298A	10634
x"00",	-- Hex Addr	298B	10635
x"00",	-- Hex Addr	298C	10636
x"00",	-- Hex Addr	298D	10637
x"00",	-- Hex Addr	298E	10638
x"00",	-- Hex Addr	298F	10639
x"00",	-- Hex Addr	2990	10640
x"00",	-- Hex Addr	2991	10641
x"00",	-- Hex Addr	2992	10642
x"00",	-- Hex Addr	2993	10643
x"00",	-- Hex Addr	2994	10644
x"00",	-- Hex Addr	2995	10645
x"00",	-- Hex Addr	2996	10646
x"00",	-- Hex Addr	2997	10647
x"00",	-- Hex Addr	2998	10648
x"00",	-- Hex Addr	2999	10649
x"00",	-- Hex Addr	299A	10650
x"00",	-- Hex Addr	299B	10651
x"00",	-- Hex Addr	299C	10652
x"00",	-- Hex Addr	299D	10653
x"00",	-- Hex Addr	299E	10654
x"00",	-- Hex Addr	299F	10655
x"00",	-- Hex Addr	29A0	10656
x"00",	-- Hex Addr	29A1	10657
x"00",	-- Hex Addr	29A2	10658
x"00",	-- Hex Addr	29A3	10659
x"00",	-- Hex Addr	29A4	10660
x"00",	-- Hex Addr	29A5	10661
x"00",	-- Hex Addr	29A6	10662
x"00",	-- Hex Addr	29A7	10663
x"00",	-- Hex Addr	29A8	10664
x"00",	-- Hex Addr	29A9	10665
x"00",	-- Hex Addr	29AA	10666
x"00",	-- Hex Addr	29AB	10667
x"00",	-- Hex Addr	29AC	10668
x"00",	-- Hex Addr	29AD	10669
x"00",	-- Hex Addr	29AE	10670
x"00",	-- Hex Addr	29AF	10671
x"00",	-- Hex Addr	29B0	10672
x"00",	-- Hex Addr	29B1	10673
x"00",	-- Hex Addr	29B2	10674
x"00",	-- Hex Addr	29B3	10675
x"00",	-- Hex Addr	29B4	10676
x"00",	-- Hex Addr	29B5	10677
x"00",	-- Hex Addr	29B6	10678
x"00",	-- Hex Addr	29B7	10679
x"00",	-- Hex Addr	29B8	10680
x"00",	-- Hex Addr	29B9	10681
x"00",	-- Hex Addr	29BA	10682
x"00",	-- Hex Addr	29BB	10683
x"00",	-- Hex Addr	29BC	10684
x"00",	-- Hex Addr	29BD	10685
x"00",	-- Hex Addr	29BE	10686
x"00",	-- Hex Addr	29BF	10687
x"00",	-- Hex Addr	29C0	10688
x"00",	-- Hex Addr	29C1	10689
x"00",	-- Hex Addr	29C2	10690
x"00",	-- Hex Addr	29C3	10691
x"00",	-- Hex Addr	29C4	10692
x"00",	-- Hex Addr	29C5	10693
x"00",	-- Hex Addr	29C6	10694
x"00",	-- Hex Addr	29C7	10695
x"00",	-- Hex Addr	29C8	10696
x"00",	-- Hex Addr	29C9	10697
x"00",	-- Hex Addr	29CA	10698
x"00",	-- Hex Addr	29CB	10699
x"00",	-- Hex Addr	29CC	10700
x"00",	-- Hex Addr	29CD	10701
x"00",	-- Hex Addr	29CE	10702
x"00",	-- Hex Addr	29CF	10703
x"00",	-- Hex Addr	29D0	10704
x"00",	-- Hex Addr	29D1	10705
x"00",	-- Hex Addr	29D2	10706
x"00",	-- Hex Addr	29D3	10707
x"00",	-- Hex Addr	29D4	10708
x"00",	-- Hex Addr	29D5	10709
x"00",	-- Hex Addr	29D6	10710
x"00",	-- Hex Addr	29D7	10711
x"00",	-- Hex Addr	29D8	10712
x"00",	-- Hex Addr	29D9	10713
x"00",	-- Hex Addr	29DA	10714
x"00",	-- Hex Addr	29DB	10715
x"00",	-- Hex Addr	29DC	10716
x"00",	-- Hex Addr	29DD	10717
x"00",	-- Hex Addr	29DE	10718
x"00",	-- Hex Addr	29DF	10719
x"00",	-- Hex Addr	29E0	10720
x"00",	-- Hex Addr	29E1	10721
x"00",	-- Hex Addr	29E2	10722
x"00",	-- Hex Addr	29E3	10723
x"00",	-- Hex Addr	29E4	10724
x"00",	-- Hex Addr	29E5	10725
x"00",	-- Hex Addr	29E6	10726
x"00",	-- Hex Addr	29E7	10727
x"00",	-- Hex Addr	29E8	10728
x"00",	-- Hex Addr	29E9	10729
x"00",	-- Hex Addr	29EA	10730
x"00",	-- Hex Addr	29EB	10731
x"00",	-- Hex Addr	29EC	10732
x"00",	-- Hex Addr	29ED	10733
x"00",	-- Hex Addr	29EE	10734
x"00",	-- Hex Addr	29EF	10735
x"00",	-- Hex Addr	29F0	10736
x"00",	-- Hex Addr	29F1	10737
x"00",	-- Hex Addr	29F2	10738
x"00",	-- Hex Addr	29F3	10739
x"00",	-- Hex Addr	29F4	10740
x"00",	-- Hex Addr	29F5	10741
x"00",	-- Hex Addr	29F6	10742
x"00",	-- Hex Addr	29F7	10743
x"00",	-- Hex Addr	29F8	10744
x"00",	-- Hex Addr	29F9	10745
x"00",	-- Hex Addr	29FA	10746
x"00",	-- Hex Addr	29FB	10747
x"00",	-- Hex Addr	29FC	10748
x"00",	-- Hex Addr	29FD	10749
x"00",	-- Hex Addr	29FE	10750
x"00",	-- Hex Addr	29FF	10751
x"00",	-- Hex Addr	2A00	10752
x"00",	-- Hex Addr	2A01	10753
x"00",	-- Hex Addr	2A02	10754
x"00",	-- Hex Addr	2A03	10755
x"00",	-- Hex Addr	2A04	10756
x"00",	-- Hex Addr	2A05	10757
x"00",	-- Hex Addr	2A06	10758
x"00",	-- Hex Addr	2A07	10759
x"00",	-- Hex Addr	2A08	10760
x"00",	-- Hex Addr	2A09	10761
x"00",	-- Hex Addr	2A0A	10762
x"00",	-- Hex Addr	2A0B	10763
x"00",	-- Hex Addr	2A0C	10764
x"00",	-- Hex Addr	2A0D	10765
x"00",	-- Hex Addr	2A0E	10766
x"00",	-- Hex Addr	2A0F	10767
x"00",	-- Hex Addr	2A10	10768
x"00",	-- Hex Addr	2A11	10769
x"00",	-- Hex Addr	2A12	10770
x"00",	-- Hex Addr	2A13	10771
x"00",	-- Hex Addr	2A14	10772
x"00",	-- Hex Addr	2A15	10773
x"00",	-- Hex Addr	2A16	10774
x"00",	-- Hex Addr	2A17	10775
x"00",	-- Hex Addr	2A18	10776
x"00",	-- Hex Addr	2A19	10777
x"00",	-- Hex Addr	2A1A	10778
x"00",	-- Hex Addr	2A1B	10779
x"00",	-- Hex Addr	2A1C	10780
x"00",	-- Hex Addr	2A1D	10781
x"00",	-- Hex Addr	2A1E	10782
x"00",	-- Hex Addr	2A1F	10783
x"00",	-- Hex Addr	2A20	10784
x"00",	-- Hex Addr	2A21	10785
x"00",	-- Hex Addr	2A22	10786
x"00",	-- Hex Addr	2A23	10787
x"00",	-- Hex Addr	2A24	10788
x"00",	-- Hex Addr	2A25	10789
x"00",	-- Hex Addr	2A26	10790
x"00",	-- Hex Addr	2A27	10791
x"00",	-- Hex Addr	2A28	10792
x"00",	-- Hex Addr	2A29	10793
x"00",	-- Hex Addr	2A2A	10794
x"00",	-- Hex Addr	2A2B	10795
x"00",	-- Hex Addr	2A2C	10796
x"00",	-- Hex Addr	2A2D	10797
x"00",	-- Hex Addr	2A2E	10798
x"00",	-- Hex Addr	2A2F	10799
x"00",	-- Hex Addr	2A30	10800
x"00",	-- Hex Addr	2A31	10801
x"00",	-- Hex Addr	2A32	10802
x"00",	-- Hex Addr	2A33	10803
x"00",	-- Hex Addr	2A34	10804
x"00",	-- Hex Addr	2A35	10805
x"00",	-- Hex Addr	2A36	10806
x"00",	-- Hex Addr	2A37	10807
x"00",	-- Hex Addr	2A38	10808
x"00",	-- Hex Addr	2A39	10809
x"00",	-- Hex Addr	2A3A	10810
x"00",	-- Hex Addr	2A3B	10811
x"00",	-- Hex Addr	2A3C	10812
x"00",	-- Hex Addr	2A3D	10813
x"00",	-- Hex Addr	2A3E	10814
x"00",	-- Hex Addr	2A3F	10815
x"00",	-- Hex Addr	2A40	10816
x"00",	-- Hex Addr	2A41	10817
x"00",	-- Hex Addr	2A42	10818
x"00",	-- Hex Addr	2A43	10819
x"00",	-- Hex Addr	2A44	10820
x"00",	-- Hex Addr	2A45	10821
x"00",	-- Hex Addr	2A46	10822
x"00",	-- Hex Addr	2A47	10823
x"00",	-- Hex Addr	2A48	10824
x"00",	-- Hex Addr	2A49	10825
x"00",	-- Hex Addr	2A4A	10826
x"00",	-- Hex Addr	2A4B	10827
x"00",	-- Hex Addr	2A4C	10828
x"00",	-- Hex Addr	2A4D	10829
x"00",	-- Hex Addr	2A4E	10830
x"00",	-- Hex Addr	2A4F	10831
x"00",	-- Hex Addr	2A50	10832
x"00",	-- Hex Addr	2A51	10833
x"00",	-- Hex Addr	2A52	10834
x"00",	-- Hex Addr	2A53	10835
x"00",	-- Hex Addr	2A54	10836
x"00",	-- Hex Addr	2A55	10837
x"00",	-- Hex Addr	2A56	10838
x"00",	-- Hex Addr	2A57	10839
x"00",	-- Hex Addr	2A58	10840
x"00",	-- Hex Addr	2A59	10841
x"00",	-- Hex Addr	2A5A	10842
x"00",	-- Hex Addr	2A5B	10843
x"00",	-- Hex Addr	2A5C	10844
x"00",	-- Hex Addr	2A5D	10845
x"00",	-- Hex Addr	2A5E	10846
x"00",	-- Hex Addr	2A5F	10847
x"00",	-- Hex Addr	2A60	10848
x"00",	-- Hex Addr	2A61	10849
x"00",	-- Hex Addr	2A62	10850
x"00",	-- Hex Addr	2A63	10851
x"00",	-- Hex Addr	2A64	10852
x"00",	-- Hex Addr	2A65	10853
x"00",	-- Hex Addr	2A66	10854
x"00",	-- Hex Addr	2A67	10855
x"00",	-- Hex Addr	2A68	10856
x"00",	-- Hex Addr	2A69	10857
x"00",	-- Hex Addr	2A6A	10858
x"00",	-- Hex Addr	2A6B	10859
x"00",	-- Hex Addr	2A6C	10860
x"00",	-- Hex Addr	2A6D	10861
x"00",	-- Hex Addr	2A6E	10862
x"00",	-- Hex Addr	2A6F	10863
x"00",	-- Hex Addr	2A70	10864
x"00",	-- Hex Addr	2A71	10865
x"00",	-- Hex Addr	2A72	10866
x"00",	-- Hex Addr	2A73	10867
x"00",	-- Hex Addr	2A74	10868
x"00",	-- Hex Addr	2A75	10869
x"00",	-- Hex Addr	2A76	10870
x"00",	-- Hex Addr	2A77	10871
x"00",	-- Hex Addr	2A78	10872
x"00",	-- Hex Addr	2A79	10873
x"00",	-- Hex Addr	2A7A	10874
x"00",	-- Hex Addr	2A7B	10875
x"00",	-- Hex Addr	2A7C	10876
x"00",	-- Hex Addr	2A7D	10877
x"00",	-- Hex Addr	2A7E	10878
x"00",	-- Hex Addr	2A7F	10879
x"00",	-- Hex Addr	2A80	10880
x"00",	-- Hex Addr	2A81	10881
x"00",	-- Hex Addr	2A82	10882
x"00",	-- Hex Addr	2A83	10883
x"00",	-- Hex Addr	2A84	10884
x"00",	-- Hex Addr	2A85	10885
x"00",	-- Hex Addr	2A86	10886
x"00",	-- Hex Addr	2A87	10887
x"00",	-- Hex Addr	2A88	10888
x"00",	-- Hex Addr	2A89	10889
x"00",	-- Hex Addr	2A8A	10890
x"00",	-- Hex Addr	2A8B	10891
x"00",	-- Hex Addr	2A8C	10892
x"00",	-- Hex Addr	2A8D	10893
x"00",	-- Hex Addr	2A8E	10894
x"00",	-- Hex Addr	2A8F	10895
x"00",	-- Hex Addr	2A90	10896
x"00",	-- Hex Addr	2A91	10897
x"00",	-- Hex Addr	2A92	10898
x"00",	-- Hex Addr	2A93	10899
x"00",	-- Hex Addr	2A94	10900
x"00",	-- Hex Addr	2A95	10901
x"00",	-- Hex Addr	2A96	10902
x"00",	-- Hex Addr	2A97	10903
x"00",	-- Hex Addr	2A98	10904
x"00",	-- Hex Addr	2A99	10905
x"00",	-- Hex Addr	2A9A	10906
x"00",	-- Hex Addr	2A9B	10907
x"00",	-- Hex Addr	2A9C	10908
x"00",	-- Hex Addr	2A9D	10909
x"00",	-- Hex Addr	2A9E	10910
x"00",	-- Hex Addr	2A9F	10911
x"00",	-- Hex Addr	2AA0	10912
x"00",	-- Hex Addr	2AA1	10913
x"00",	-- Hex Addr	2AA2	10914
x"00",	-- Hex Addr	2AA3	10915
x"00",	-- Hex Addr	2AA4	10916
x"00",	-- Hex Addr	2AA5	10917
x"00",	-- Hex Addr	2AA6	10918
x"00",	-- Hex Addr	2AA7	10919
x"00",	-- Hex Addr	2AA8	10920
x"00",	-- Hex Addr	2AA9	10921
x"00",	-- Hex Addr	2AAA	10922
x"00",	-- Hex Addr	2AAB	10923
x"00",	-- Hex Addr	2AAC	10924
x"00",	-- Hex Addr	2AAD	10925
x"00",	-- Hex Addr	2AAE	10926
x"00",	-- Hex Addr	2AAF	10927
x"00",	-- Hex Addr	2AB0	10928
x"00",	-- Hex Addr	2AB1	10929
x"00",	-- Hex Addr	2AB2	10930
x"00",	-- Hex Addr	2AB3	10931
x"00",	-- Hex Addr	2AB4	10932
x"00",	-- Hex Addr	2AB5	10933
x"00",	-- Hex Addr	2AB6	10934
x"00",	-- Hex Addr	2AB7	10935
x"00",	-- Hex Addr	2AB8	10936
x"00",	-- Hex Addr	2AB9	10937
x"00",	-- Hex Addr	2ABA	10938
x"00",	-- Hex Addr	2ABB	10939
x"00",	-- Hex Addr	2ABC	10940
x"00",	-- Hex Addr	2ABD	10941
x"00",	-- Hex Addr	2ABE	10942
x"00",	-- Hex Addr	2ABF	10943
x"00",	-- Hex Addr	2AC0	10944
x"00",	-- Hex Addr	2AC1	10945
x"00",	-- Hex Addr	2AC2	10946
x"00",	-- Hex Addr	2AC3	10947
x"00",	-- Hex Addr	2AC4	10948
x"00",	-- Hex Addr	2AC5	10949
x"00",	-- Hex Addr	2AC6	10950
x"00",	-- Hex Addr	2AC7	10951
x"00",	-- Hex Addr	2AC8	10952
x"00",	-- Hex Addr	2AC9	10953
x"00",	-- Hex Addr	2ACA	10954
x"00",	-- Hex Addr	2ACB	10955
x"00",	-- Hex Addr	2ACC	10956
x"00",	-- Hex Addr	2ACD	10957
x"00",	-- Hex Addr	2ACE	10958
x"00",	-- Hex Addr	2ACF	10959
x"00",	-- Hex Addr	2AD0	10960
x"00",	-- Hex Addr	2AD1	10961
x"00",	-- Hex Addr	2AD2	10962
x"00",	-- Hex Addr	2AD3	10963
x"00",	-- Hex Addr	2AD4	10964
x"00",	-- Hex Addr	2AD5	10965
x"00",	-- Hex Addr	2AD6	10966
x"00",	-- Hex Addr	2AD7	10967
x"00",	-- Hex Addr	2AD8	10968
x"00",	-- Hex Addr	2AD9	10969
x"00",	-- Hex Addr	2ADA	10970
x"00",	-- Hex Addr	2ADB	10971
x"00",	-- Hex Addr	2ADC	10972
x"00",	-- Hex Addr	2ADD	10973
x"00",	-- Hex Addr	2ADE	10974
x"00",	-- Hex Addr	2ADF	10975
x"00",	-- Hex Addr	2AE0	10976
x"00",	-- Hex Addr	2AE1	10977
x"00",	-- Hex Addr	2AE2	10978
x"00",	-- Hex Addr	2AE3	10979
x"00",	-- Hex Addr	2AE4	10980
x"00",	-- Hex Addr	2AE5	10981
x"00",	-- Hex Addr	2AE6	10982
x"00",	-- Hex Addr	2AE7	10983
x"00",	-- Hex Addr	2AE8	10984
x"00",	-- Hex Addr	2AE9	10985
x"00",	-- Hex Addr	2AEA	10986
x"00",	-- Hex Addr	2AEB	10987
x"00",	-- Hex Addr	2AEC	10988
x"00",	-- Hex Addr	2AED	10989
x"00",	-- Hex Addr	2AEE	10990
x"00",	-- Hex Addr	2AEF	10991
x"00",	-- Hex Addr	2AF0	10992
x"00",	-- Hex Addr	2AF1	10993
x"00",	-- Hex Addr	2AF2	10994
x"00",	-- Hex Addr	2AF3	10995
x"00",	-- Hex Addr	2AF4	10996
x"00",	-- Hex Addr	2AF5	10997
x"00",	-- Hex Addr	2AF6	10998
x"00",	-- Hex Addr	2AF7	10999
x"00",	-- Hex Addr	2AF8	11000
x"00",	-- Hex Addr	2AF9	11001
x"00",	-- Hex Addr	2AFA	11002
x"00",	-- Hex Addr	2AFB	11003
x"00",	-- Hex Addr	2AFC	11004
x"00",	-- Hex Addr	2AFD	11005
x"00",	-- Hex Addr	2AFE	11006
x"00",	-- Hex Addr	2AFF	11007
x"00",	-- Hex Addr	2B00	11008
x"00",	-- Hex Addr	2B01	11009
x"00",	-- Hex Addr	2B02	11010
x"00",	-- Hex Addr	2B03	11011
x"00",	-- Hex Addr	2B04	11012
x"00",	-- Hex Addr	2B05	11013
x"00",	-- Hex Addr	2B06	11014
x"00",	-- Hex Addr	2B07	11015
x"00",	-- Hex Addr	2B08	11016
x"00",	-- Hex Addr	2B09	11017
x"00",	-- Hex Addr	2B0A	11018
x"00",	-- Hex Addr	2B0B	11019
x"00",	-- Hex Addr	2B0C	11020
x"00",	-- Hex Addr	2B0D	11021
x"00",	-- Hex Addr	2B0E	11022
x"00",	-- Hex Addr	2B0F	11023
x"00",	-- Hex Addr	2B10	11024
x"00",	-- Hex Addr	2B11	11025
x"00",	-- Hex Addr	2B12	11026
x"00",	-- Hex Addr	2B13	11027
x"00",	-- Hex Addr	2B14	11028
x"00",	-- Hex Addr	2B15	11029
x"00",	-- Hex Addr	2B16	11030
x"00",	-- Hex Addr	2B17	11031
x"00",	-- Hex Addr	2B18	11032
x"00",	-- Hex Addr	2B19	11033
x"00",	-- Hex Addr	2B1A	11034
x"00",	-- Hex Addr	2B1B	11035
x"00",	-- Hex Addr	2B1C	11036
x"00",	-- Hex Addr	2B1D	11037
x"00",	-- Hex Addr	2B1E	11038
x"00",	-- Hex Addr	2B1F	11039
x"00",	-- Hex Addr	2B20	11040
x"00",	-- Hex Addr	2B21	11041
x"00",	-- Hex Addr	2B22	11042
x"00",	-- Hex Addr	2B23	11043
x"00",	-- Hex Addr	2B24	11044
x"00",	-- Hex Addr	2B25	11045
x"00",	-- Hex Addr	2B26	11046
x"00",	-- Hex Addr	2B27	11047
x"00",	-- Hex Addr	2B28	11048
x"00",	-- Hex Addr	2B29	11049
x"00",	-- Hex Addr	2B2A	11050
x"00",	-- Hex Addr	2B2B	11051
x"00",	-- Hex Addr	2B2C	11052
x"00",	-- Hex Addr	2B2D	11053
x"00",	-- Hex Addr	2B2E	11054
x"00",	-- Hex Addr	2B2F	11055
x"00",	-- Hex Addr	2B30	11056
x"00",	-- Hex Addr	2B31	11057
x"00",	-- Hex Addr	2B32	11058
x"00",	-- Hex Addr	2B33	11059
x"00",	-- Hex Addr	2B34	11060
x"00",	-- Hex Addr	2B35	11061
x"00",	-- Hex Addr	2B36	11062
x"00",	-- Hex Addr	2B37	11063
x"00",	-- Hex Addr	2B38	11064
x"00",	-- Hex Addr	2B39	11065
x"00",	-- Hex Addr	2B3A	11066
x"00",	-- Hex Addr	2B3B	11067
x"00",	-- Hex Addr	2B3C	11068
x"00",	-- Hex Addr	2B3D	11069
x"00",	-- Hex Addr	2B3E	11070
x"00",	-- Hex Addr	2B3F	11071
x"00",	-- Hex Addr	2B40	11072
x"00",	-- Hex Addr	2B41	11073
x"00",	-- Hex Addr	2B42	11074
x"00",	-- Hex Addr	2B43	11075
x"00",	-- Hex Addr	2B44	11076
x"00",	-- Hex Addr	2B45	11077
x"00",	-- Hex Addr	2B46	11078
x"00",	-- Hex Addr	2B47	11079
x"00",	-- Hex Addr	2B48	11080
x"00",	-- Hex Addr	2B49	11081
x"00",	-- Hex Addr	2B4A	11082
x"00",	-- Hex Addr	2B4B	11083
x"00",	-- Hex Addr	2B4C	11084
x"00",	-- Hex Addr	2B4D	11085
x"00",	-- Hex Addr	2B4E	11086
x"00",	-- Hex Addr	2B4F	11087
x"00",	-- Hex Addr	2B50	11088
x"00",	-- Hex Addr	2B51	11089
x"00",	-- Hex Addr	2B52	11090
x"00",	-- Hex Addr	2B53	11091
x"00",	-- Hex Addr	2B54	11092
x"00",	-- Hex Addr	2B55	11093
x"00",	-- Hex Addr	2B56	11094
x"00",	-- Hex Addr	2B57	11095
x"00",	-- Hex Addr	2B58	11096
x"00",	-- Hex Addr	2B59	11097
x"00",	-- Hex Addr	2B5A	11098
x"00",	-- Hex Addr	2B5B	11099
x"00",	-- Hex Addr	2B5C	11100
x"00",	-- Hex Addr	2B5D	11101
x"00",	-- Hex Addr	2B5E	11102
x"00",	-- Hex Addr	2B5F	11103
x"00",	-- Hex Addr	2B60	11104
x"00",	-- Hex Addr	2B61	11105
x"00",	-- Hex Addr	2B62	11106
x"00",	-- Hex Addr	2B63	11107
x"00",	-- Hex Addr	2B64	11108
x"00",	-- Hex Addr	2B65	11109
x"00",	-- Hex Addr	2B66	11110
x"00",	-- Hex Addr	2B67	11111
x"00",	-- Hex Addr	2B68	11112
x"00",	-- Hex Addr	2B69	11113
x"00",	-- Hex Addr	2B6A	11114
x"00",	-- Hex Addr	2B6B	11115
x"00",	-- Hex Addr	2B6C	11116
x"00",	-- Hex Addr	2B6D	11117
x"00",	-- Hex Addr	2B6E	11118
x"00",	-- Hex Addr	2B6F	11119
x"00",	-- Hex Addr	2B70	11120
x"00",	-- Hex Addr	2B71	11121
x"00",	-- Hex Addr	2B72	11122
x"00",	-- Hex Addr	2B73	11123
x"00",	-- Hex Addr	2B74	11124
x"00",	-- Hex Addr	2B75	11125
x"00",	-- Hex Addr	2B76	11126
x"00",	-- Hex Addr	2B77	11127
x"00",	-- Hex Addr	2B78	11128
x"00",	-- Hex Addr	2B79	11129
x"00",	-- Hex Addr	2B7A	11130
x"00",	-- Hex Addr	2B7B	11131
x"00",	-- Hex Addr	2B7C	11132
x"00",	-- Hex Addr	2B7D	11133
x"00",	-- Hex Addr	2B7E	11134
x"00",	-- Hex Addr	2B7F	11135
x"00",	-- Hex Addr	2B80	11136
x"00",	-- Hex Addr	2B81	11137
x"00",	-- Hex Addr	2B82	11138
x"00",	-- Hex Addr	2B83	11139
x"00",	-- Hex Addr	2B84	11140
x"00",	-- Hex Addr	2B85	11141
x"00",	-- Hex Addr	2B86	11142
x"00",	-- Hex Addr	2B87	11143
x"00",	-- Hex Addr	2B88	11144
x"00",	-- Hex Addr	2B89	11145
x"00",	-- Hex Addr	2B8A	11146
x"00",	-- Hex Addr	2B8B	11147
x"00",	-- Hex Addr	2B8C	11148
x"00",	-- Hex Addr	2B8D	11149
x"00",	-- Hex Addr	2B8E	11150
x"00",	-- Hex Addr	2B8F	11151
x"00",	-- Hex Addr	2B90	11152
x"00",	-- Hex Addr	2B91	11153
x"00",	-- Hex Addr	2B92	11154
x"00",	-- Hex Addr	2B93	11155
x"00",	-- Hex Addr	2B94	11156
x"00",	-- Hex Addr	2B95	11157
x"00",	-- Hex Addr	2B96	11158
x"00",	-- Hex Addr	2B97	11159
x"00",	-- Hex Addr	2B98	11160
x"00",	-- Hex Addr	2B99	11161
x"00",	-- Hex Addr	2B9A	11162
x"00",	-- Hex Addr	2B9B	11163
x"00",	-- Hex Addr	2B9C	11164
x"00",	-- Hex Addr	2B9D	11165
x"00",	-- Hex Addr	2B9E	11166
x"00",	-- Hex Addr	2B9F	11167
x"00",	-- Hex Addr	2BA0	11168
x"00",	-- Hex Addr	2BA1	11169
x"00",	-- Hex Addr	2BA2	11170
x"00",	-- Hex Addr	2BA3	11171
x"00",	-- Hex Addr	2BA4	11172
x"00",	-- Hex Addr	2BA5	11173
x"00",	-- Hex Addr	2BA6	11174
x"00",	-- Hex Addr	2BA7	11175
x"00",	-- Hex Addr	2BA8	11176
x"00",	-- Hex Addr	2BA9	11177
x"00",	-- Hex Addr	2BAA	11178
x"00",	-- Hex Addr	2BAB	11179
x"00",	-- Hex Addr	2BAC	11180
x"00",	-- Hex Addr	2BAD	11181
x"00",	-- Hex Addr	2BAE	11182
x"00",	-- Hex Addr	2BAF	11183
x"00",	-- Hex Addr	2BB0	11184
x"00",	-- Hex Addr	2BB1	11185
x"00",	-- Hex Addr	2BB2	11186
x"00",	-- Hex Addr	2BB3	11187
x"00",	-- Hex Addr	2BB4	11188
x"00",	-- Hex Addr	2BB5	11189
x"00",	-- Hex Addr	2BB6	11190
x"00",	-- Hex Addr	2BB7	11191
x"00",	-- Hex Addr	2BB8	11192
x"00",	-- Hex Addr	2BB9	11193
x"00",	-- Hex Addr	2BBA	11194
x"00",	-- Hex Addr	2BBB	11195
x"00",	-- Hex Addr	2BBC	11196
x"00",	-- Hex Addr	2BBD	11197
x"00",	-- Hex Addr	2BBE	11198
x"00",	-- Hex Addr	2BBF	11199
x"00",	-- Hex Addr	2BC0	11200
x"00",	-- Hex Addr	2BC1	11201
x"00",	-- Hex Addr	2BC2	11202
x"00",	-- Hex Addr	2BC3	11203
x"00",	-- Hex Addr	2BC4	11204
x"00",	-- Hex Addr	2BC5	11205
x"00",	-- Hex Addr	2BC6	11206
x"00",	-- Hex Addr	2BC7	11207
x"00",	-- Hex Addr	2BC8	11208
x"00",	-- Hex Addr	2BC9	11209
x"00",	-- Hex Addr	2BCA	11210
x"00",	-- Hex Addr	2BCB	11211
x"00",	-- Hex Addr	2BCC	11212
x"00",	-- Hex Addr	2BCD	11213
x"00",	-- Hex Addr	2BCE	11214
x"00",	-- Hex Addr	2BCF	11215
x"00",	-- Hex Addr	2BD0	11216
x"00",	-- Hex Addr	2BD1	11217
x"00",	-- Hex Addr	2BD2	11218
x"00",	-- Hex Addr	2BD3	11219
x"00",	-- Hex Addr	2BD4	11220
x"00",	-- Hex Addr	2BD5	11221
x"00",	-- Hex Addr	2BD6	11222
x"00",	-- Hex Addr	2BD7	11223
x"00",	-- Hex Addr	2BD8	11224
x"00",	-- Hex Addr	2BD9	11225
x"00",	-- Hex Addr	2BDA	11226
x"00",	-- Hex Addr	2BDB	11227
x"00",	-- Hex Addr	2BDC	11228
x"00",	-- Hex Addr	2BDD	11229
x"00",	-- Hex Addr	2BDE	11230
x"00",	-- Hex Addr	2BDF	11231
x"00",	-- Hex Addr	2BE0	11232
x"00",	-- Hex Addr	2BE1	11233
x"00",	-- Hex Addr	2BE2	11234
x"00",	-- Hex Addr	2BE3	11235
x"00",	-- Hex Addr	2BE4	11236
x"00",	-- Hex Addr	2BE5	11237
x"00",	-- Hex Addr	2BE6	11238
x"00",	-- Hex Addr	2BE7	11239
x"00",	-- Hex Addr	2BE8	11240
x"00",	-- Hex Addr	2BE9	11241
x"00",	-- Hex Addr	2BEA	11242
x"00",	-- Hex Addr	2BEB	11243
x"00",	-- Hex Addr	2BEC	11244
x"00",	-- Hex Addr	2BED	11245
x"00",	-- Hex Addr	2BEE	11246
x"00",	-- Hex Addr	2BEF	11247
x"00",	-- Hex Addr	2BF0	11248
x"00",	-- Hex Addr	2BF1	11249
x"00",	-- Hex Addr	2BF2	11250
x"00",	-- Hex Addr	2BF3	11251
x"00",	-- Hex Addr	2BF4	11252
x"00",	-- Hex Addr	2BF5	11253
x"00",	-- Hex Addr	2BF6	11254
x"00",	-- Hex Addr	2BF7	11255
x"00",	-- Hex Addr	2BF8	11256
x"00",	-- Hex Addr	2BF9	11257
x"00",	-- Hex Addr	2BFA	11258
x"00",	-- Hex Addr	2BFB	11259
x"00",	-- Hex Addr	2BFC	11260
x"00",	-- Hex Addr	2BFD	11261
x"00",	-- Hex Addr	2BFE	11262
x"00",	-- Hex Addr	2BFF	11263
x"00",	-- Hex Addr	2C00	11264
x"00",	-- Hex Addr	2C01	11265
x"00",	-- Hex Addr	2C02	11266
x"00",	-- Hex Addr	2C03	11267
x"00",	-- Hex Addr	2C04	11268
x"00",	-- Hex Addr	2C05	11269
x"00",	-- Hex Addr	2C06	11270
x"00",	-- Hex Addr	2C07	11271
x"00",	-- Hex Addr	2C08	11272
x"00",	-- Hex Addr	2C09	11273
x"00",	-- Hex Addr	2C0A	11274
x"00",	-- Hex Addr	2C0B	11275
x"00",	-- Hex Addr	2C0C	11276
x"00",	-- Hex Addr	2C0D	11277
x"00",	-- Hex Addr	2C0E	11278
x"00",	-- Hex Addr	2C0F	11279
x"00",	-- Hex Addr	2C10	11280
x"00",	-- Hex Addr	2C11	11281
x"00",	-- Hex Addr	2C12	11282
x"00",	-- Hex Addr	2C13	11283
x"00",	-- Hex Addr	2C14	11284
x"00",	-- Hex Addr	2C15	11285
x"00",	-- Hex Addr	2C16	11286
x"00",	-- Hex Addr	2C17	11287
x"00",	-- Hex Addr	2C18	11288
x"00",	-- Hex Addr	2C19	11289
x"00",	-- Hex Addr	2C1A	11290
x"00",	-- Hex Addr	2C1B	11291
x"00",	-- Hex Addr	2C1C	11292
x"00",	-- Hex Addr	2C1D	11293
x"00",	-- Hex Addr	2C1E	11294
x"00",	-- Hex Addr	2C1F	11295
x"00",	-- Hex Addr	2C20	11296
x"00",	-- Hex Addr	2C21	11297
x"00",	-- Hex Addr	2C22	11298
x"00",	-- Hex Addr	2C23	11299
x"00",	-- Hex Addr	2C24	11300
x"00",	-- Hex Addr	2C25	11301
x"00",	-- Hex Addr	2C26	11302
x"00",	-- Hex Addr	2C27	11303
x"00",	-- Hex Addr	2C28	11304
x"00",	-- Hex Addr	2C29	11305
x"00",	-- Hex Addr	2C2A	11306
x"00",	-- Hex Addr	2C2B	11307
x"00",	-- Hex Addr	2C2C	11308
x"00",	-- Hex Addr	2C2D	11309
x"00",	-- Hex Addr	2C2E	11310
x"00",	-- Hex Addr	2C2F	11311
x"00",	-- Hex Addr	2C30	11312
x"00",	-- Hex Addr	2C31	11313
x"00",	-- Hex Addr	2C32	11314
x"00",	-- Hex Addr	2C33	11315
x"00",	-- Hex Addr	2C34	11316
x"00",	-- Hex Addr	2C35	11317
x"00",	-- Hex Addr	2C36	11318
x"00",	-- Hex Addr	2C37	11319
x"00",	-- Hex Addr	2C38	11320
x"00",	-- Hex Addr	2C39	11321
x"00",	-- Hex Addr	2C3A	11322
x"00",	-- Hex Addr	2C3B	11323
x"00",	-- Hex Addr	2C3C	11324
x"00",	-- Hex Addr	2C3D	11325
x"00",	-- Hex Addr	2C3E	11326
x"00",	-- Hex Addr	2C3F	11327
x"00",	-- Hex Addr	2C40	11328
x"00",	-- Hex Addr	2C41	11329
x"00",	-- Hex Addr	2C42	11330
x"00",	-- Hex Addr	2C43	11331
x"00",	-- Hex Addr	2C44	11332
x"00",	-- Hex Addr	2C45	11333
x"00",	-- Hex Addr	2C46	11334
x"00",	-- Hex Addr	2C47	11335
x"00",	-- Hex Addr	2C48	11336
x"00",	-- Hex Addr	2C49	11337
x"00",	-- Hex Addr	2C4A	11338
x"00",	-- Hex Addr	2C4B	11339
x"00",	-- Hex Addr	2C4C	11340
x"00",	-- Hex Addr	2C4D	11341
x"00",	-- Hex Addr	2C4E	11342
x"00",	-- Hex Addr	2C4F	11343
x"00",	-- Hex Addr	2C50	11344
x"00",	-- Hex Addr	2C51	11345
x"00",	-- Hex Addr	2C52	11346
x"00",	-- Hex Addr	2C53	11347
x"00",	-- Hex Addr	2C54	11348
x"00",	-- Hex Addr	2C55	11349
x"00",	-- Hex Addr	2C56	11350
x"00",	-- Hex Addr	2C57	11351
x"00",	-- Hex Addr	2C58	11352
x"00",	-- Hex Addr	2C59	11353
x"00",	-- Hex Addr	2C5A	11354
x"00",	-- Hex Addr	2C5B	11355
x"00",	-- Hex Addr	2C5C	11356
x"00",	-- Hex Addr	2C5D	11357
x"00",	-- Hex Addr	2C5E	11358
x"00",	-- Hex Addr	2C5F	11359
x"00",	-- Hex Addr	2C60	11360
x"00",	-- Hex Addr	2C61	11361
x"00",	-- Hex Addr	2C62	11362
x"00",	-- Hex Addr	2C63	11363
x"00",	-- Hex Addr	2C64	11364
x"00",	-- Hex Addr	2C65	11365
x"00",	-- Hex Addr	2C66	11366
x"00",	-- Hex Addr	2C67	11367
x"00",	-- Hex Addr	2C68	11368
x"00",	-- Hex Addr	2C69	11369
x"00",	-- Hex Addr	2C6A	11370
x"00",	-- Hex Addr	2C6B	11371
x"00",	-- Hex Addr	2C6C	11372
x"00",	-- Hex Addr	2C6D	11373
x"00",	-- Hex Addr	2C6E	11374
x"00",	-- Hex Addr	2C6F	11375
x"00",	-- Hex Addr	2C70	11376
x"00",	-- Hex Addr	2C71	11377
x"00",	-- Hex Addr	2C72	11378
x"00",	-- Hex Addr	2C73	11379
x"00",	-- Hex Addr	2C74	11380
x"00",	-- Hex Addr	2C75	11381
x"00",	-- Hex Addr	2C76	11382
x"00",	-- Hex Addr	2C77	11383
x"00",	-- Hex Addr	2C78	11384
x"00",	-- Hex Addr	2C79	11385
x"00",	-- Hex Addr	2C7A	11386
x"00",	-- Hex Addr	2C7B	11387
x"00",	-- Hex Addr	2C7C	11388
x"00",	-- Hex Addr	2C7D	11389
x"00",	-- Hex Addr	2C7E	11390
x"00",	-- Hex Addr	2C7F	11391
x"00",	-- Hex Addr	2C80	11392
x"00",	-- Hex Addr	2C81	11393
x"00",	-- Hex Addr	2C82	11394
x"00",	-- Hex Addr	2C83	11395
x"00",	-- Hex Addr	2C84	11396
x"00",	-- Hex Addr	2C85	11397
x"00",	-- Hex Addr	2C86	11398
x"00",	-- Hex Addr	2C87	11399
x"00",	-- Hex Addr	2C88	11400
x"00",	-- Hex Addr	2C89	11401
x"00",	-- Hex Addr	2C8A	11402
x"00",	-- Hex Addr	2C8B	11403
x"00",	-- Hex Addr	2C8C	11404
x"00",	-- Hex Addr	2C8D	11405
x"00",	-- Hex Addr	2C8E	11406
x"00",	-- Hex Addr	2C8F	11407
x"00",	-- Hex Addr	2C90	11408
x"00",	-- Hex Addr	2C91	11409
x"00",	-- Hex Addr	2C92	11410
x"00",	-- Hex Addr	2C93	11411
x"00",	-- Hex Addr	2C94	11412
x"00",	-- Hex Addr	2C95	11413
x"00",	-- Hex Addr	2C96	11414
x"00",	-- Hex Addr	2C97	11415
x"00",	-- Hex Addr	2C98	11416
x"00",	-- Hex Addr	2C99	11417
x"00",	-- Hex Addr	2C9A	11418
x"00",	-- Hex Addr	2C9B	11419
x"00",	-- Hex Addr	2C9C	11420
x"00",	-- Hex Addr	2C9D	11421
x"00",	-- Hex Addr	2C9E	11422
x"00",	-- Hex Addr	2C9F	11423
x"00",	-- Hex Addr	2CA0	11424
x"00",	-- Hex Addr	2CA1	11425
x"00",	-- Hex Addr	2CA2	11426
x"00",	-- Hex Addr	2CA3	11427
x"00",	-- Hex Addr	2CA4	11428
x"00",	-- Hex Addr	2CA5	11429
x"00",	-- Hex Addr	2CA6	11430
x"00",	-- Hex Addr	2CA7	11431
x"00",	-- Hex Addr	2CA8	11432
x"00",	-- Hex Addr	2CA9	11433
x"00",	-- Hex Addr	2CAA	11434
x"00",	-- Hex Addr	2CAB	11435
x"00",	-- Hex Addr	2CAC	11436
x"00",	-- Hex Addr	2CAD	11437
x"00",	-- Hex Addr	2CAE	11438
x"00",	-- Hex Addr	2CAF	11439
x"00",	-- Hex Addr	2CB0	11440
x"00",	-- Hex Addr	2CB1	11441
x"00",	-- Hex Addr	2CB2	11442
x"00",	-- Hex Addr	2CB3	11443
x"00",	-- Hex Addr	2CB4	11444
x"00",	-- Hex Addr	2CB5	11445
x"00",	-- Hex Addr	2CB6	11446
x"00",	-- Hex Addr	2CB7	11447
x"00",	-- Hex Addr	2CB8	11448
x"00",	-- Hex Addr	2CB9	11449
x"00",	-- Hex Addr	2CBA	11450
x"00",	-- Hex Addr	2CBB	11451
x"00",	-- Hex Addr	2CBC	11452
x"00",	-- Hex Addr	2CBD	11453
x"00",	-- Hex Addr	2CBE	11454
x"00",	-- Hex Addr	2CBF	11455
x"00",	-- Hex Addr	2CC0	11456
x"00",	-- Hex Addr	2CC1	11457
x"00",	-- Hex Addr	2CC2	11458
x"00",	-- Hex Addr	2CC3	11459
x"00",	-- Hex Addr	2CC4	11460
x"00",	-- Hex Addr	2CC5	11461
x"00",	-- Hex Addr	2CC6	11462
x"00",	-- Hex Addr	2CC7	11463
x"00",	-- Hex Addr	2CC8	11464
x"00",	-- Hex Addr	2CC9	11465
x"00",	-- Hex Addr	2CCA	11466
x"00",	-- Hex Addr	2CCB	11467
x"00",	-- Hex Addr	2CCC	11468
x"00",	-- Hex Addr	2CCD	11469
x"00",	-- Hex Addr	2CCE	11470
x"00",	-- Hex Addr	2CCF	11471
x"00",	-- Hex Addr	2CD0	11472
x"00",	-- Hex Addr	2CD1	11473
x"00",	-- Hex Addr	2CD2	11474
x"00",	-- Hex Addr	2CD3	11475
x"00",	-- Hex Addr	2CD4	11476
x"00",	-- Hex Addr	2CD5	11477
x"00",	-- Hex Addr	2CD6	11478
x"00",	-- Hex Addr	2CD7	11479
x"00",	-- Hex Addr	2CD8	11480
x"00",	-- Hex Addr	2CD9	11481
x"00",	-- Hex Addr	2CDA	11482
x"00",	-- Hex Addr	2CDB	11483
x"00",	-- Hex Addr	2CDC	11484
x"00",	-- Hex Addr	2CDD	11485
x"00",	-- Hex Addr	2CDE	11486
x"00",	-- Hex Addr	2CDF	11487
x"00",	-- Hex Addr	2CE0	11488
x"00",	-- Hex Addr	2CE1	11489
x"00",	-- Hex Addr	2CE2	11490
x"00",	-- Hex Addr	2CE3	11491
x"00",	-- Hex Addr	2CE4	11492
x"00",	-- Hex Addr	2CE5	11493
x"00",	-- Hex Addr	2CE6	11494
x"00",	-- Hex Addr	2CE7	11495
x"00",	-- Hex Addr	2CE8	11496
x"00",	-- Hex Addr	2CE9	11497
x"00",	-- Hex Addr	2CEA	11498
x"00",	-- Hex Addr	2CEB	11499
x"00",	-- Hex Addr	2CEC	11500
x"00",	-- Hex Addr	2CED	11501
x"00",	-- Hex Addr	2CEE	11502
x"00",	-- Hex Addr	2CEF	11503
x"00",	-- Hex Addr	2CF0	11504
x"00",	-- Hex Addr	2CF1	11505
x"00",	-- Hex Addr	2CF2	11506
x"00",	-- Hex Addr	2CF3	11507
x"00",	-- Hex Addr	2CF4	11508
x"00",	-- Hex Addr	2CF5	11509
x"00",	-- Hex Addr	2CF6	11510
x"00",	-- Hex Addr	2CF7	11511
x"00",	-- Hex Addr	2CF8	11512
x"00",	-- Hex Addr	2CF9	11513
x"00",	-- Hex Addr	2CFA	11514
x"00",	-- Hex Addr	2CFB	11515
x"00",	-- Hex Addr	2CFC	11516
x"00",	-- Hex Addr	2CFD	11517
x"00",	-- Hex Addr	2CFE	11518
x"00",	-- Hex Addr	2CFF	11519
x"00",	-- Hex Addr	2D00	11520
x"00",	-- Hex Addr	2D01	11521
x"00",	-- Hex Addr	2D02	11522
x"00",	-- Hex Addr	2D03	11523
x"00",	-- Hex Addr	2D04	11524
x"00",	-- Hex Addr	2D05	11525
x"00",	-- Hex Addr	2D06	11526
x"00",	-- Hex Addr	2D07	11527
x"00",	-- Hex Addr	2D08	11528
x"00",	-- Hex Addr	2D09	11529
x"00",	-- Hex Addr	2D0A	11530
x"00",	-- Hex Addr	2D0B	11531
x"00",	-- Hex Addr	2D0C	11532
x"00",	-- Hex Addr	2D0D	11533
x"00",	-- Hex Addr	2D0E	11534
x"00",	-- Hex Addr	2D0F	11535
x"00",	-- Hex Addr	2D10	11536
x"00",	-- Hex Addr	2D11	11537
x"00",	-- Hex Addr	2D12	11538
x"00",	-- Hex Addr	2D13	11539
x"00",	-- Hex Addr	2D14	11540
x"00",	-- Hex Addr	2D15	11541
x"00",	-- Hex Addr	2D16	11542
x"00",	-- Hex Addr	2D17	11543
x"00",	-- Hex Addr	2D18	11544
x"00",	-- Hex Addr	2D19	11545
x"00",	-- Hex Addr	2D1A	11546
x"00",	-- Hex Addr	2D1B	11547
x"00",	-- Hex Addr	2D1C	11548
x"00",	-- Hex Addr	2D1D	11549
x"00",	-- Hex Addr	2D1E	11550
x"00",	-- Hex Addr	2D1F	11551
x"00",	-- Hex Addr	2D20	11552
x"00",	-- Hex Addr	2D21	11553
x"00",	-- Hex Addr	2D22	11554
x"00",	-- Hex Addr	2D23	11555
x"00",	-- Hex Addr	2D24	11556
x"00",	-- Hex Addr	2D25	11557
x"00",	-- Hex Addr	2D26	11558
x"00",	-- Hex Addr	2D27	11559
x"00",	-- Hex Addr	2D28	11560
x"00",	-- Hex Addr	2D29	11561
x"00",	-- Hex Addr	2D2A	11562
x"00",	-- Hex Addr	2D2B	11563
x"00",	-- Hex Addr	2D2C	11564
x"00",	-- Hex Addr	2D2D	11565
x"00",	-- Hex Addr	2D2E	11566
x"00",	-- Hex Addr	2D2F	11567
x"00",	-- Hex Addr	2D30	11568
x"00",	-- Hex Addr	2D31	11569
x"00",	-- Hex Addr	2D32	11570
x"00",	-- Hex Addr	2D33	11571
x"00",	-- Hex Addr	2D34	11572
x"00",	-- Hex Addr	2D35	11573
x"00",	-- Hex Addr	2D36	11574
x"00",	-- Hex Addr	2D37	11575
x"00",	-- Hex Addr	2D38	11576
x"00",	-- Hex Addr	2D39	11577
x"00",	-- Hex Addr	2D3A	11578
x"00",	-- Hex Addr	2D3B	11579
x"00",	-- Hex Addr	2D3C	11580
x"00",	-- Hex Addr	2D3D	11581
x"00",	-- Hex Addr	2D3E	11582
x"00",	-- Hex Addr	2D3F	11583
x"00",	-- Hex Addr	2D40	11584
x"00",	-- Hex Addr	2D41	11585
x"00",	-- Hex Addr	2D42	11586
x"00",	-- Hex Addr	2D43	11587
x"00",	-- Hex Addr	2D44	11588
x"00",	-- Hex Addr	2D45	11589
x"00",	-- Hex Addr	2D46	11590
x"00",	-- Hex Addr	2D47	11591
x"00",	-- Hex Addr	2D48	11592
x"00",	-- Hex Addr	2D49	11593
x"00",	-- Hex Addr	2D4A	11594
x"00",	-- Hex Addr	2D4B	11595
x"00",	-- Hex Addr	2D4C	11596
x"00",	-- Hex Addr	2D4D	11597
x"00",	-- Hex Addr	2D4E	11598
x"00",	-- Hex Addr	2D4F	11599
x"00",	-- Hex Addr	2D50	11600
x"00",	-- Hex Addr	2D51	11601
x"00",	-- Hex Addr	2D52	11602
x"00",	-- Hex Addr	2D53	11603
x"00",	-- Hex Addr	2D54	11604
x"00",	-- Hex Addr	2D55	11605
x"00",	-- Hex Addr	2D56	11606
x"00",	-- Hex Addr	2D57	11607
x"00",	-- Hex Addr	2D58	11608
x"00",	-- Hex Addr	2D59	11609
x"00",	-- Hex Addr	2D5A	11610
x"00",	-- Hex Addr	2D5B	11611
x"00",	-- Hex Addr	2D5C	11612
x"00",	-- Hex Addr	2D5D	11613
x"00",	-- Hex Addr	2D5E	11614
x"00",	-- Hex Addr	2D5F	11615
x"00",	-- Hex Addr	2D60	11616
x"00",	-- Hex Addr	2D61	11617
x"00",	-- Hex Addr	2D62	11618
x"00",	-- Hex Addr	2D63	11619
x"00",	-- Hex Addr	2D64	11620
x"00",	-- Hex Addr	2D65	11621
x"00",	-- Hex Addr	2D66	11622
x"00",	-- Hex Addr	2D67	11623
x"00",	-- Hex Addr	2D68	11624
x"00",	-- Hex Addr	2D69	11625
x"00",	-- Hex Addr	2D6A	11626
x"00",	-- Hex Addr	2D6B	11627
x"00",	-- Hex Addr	2D6C	11628
x"00",	-- Hex Addr	2D6D	11629
x"00",	-- Hex Addr	2D6E	11630
x"00",	-- Hex Addr	2D6F	11631
x"00",	-- Hex Addr	2D70	11632
x"00",	-- Hex Addr	2D71	11633
x"00",	-- Hex Addr	2D72	11634
x"00",	-- Hex Addr	2D73	11635
x"00",	-- Hex Addr	2D74	11636
x"00",	-- Hex Addr	2D75	11637
x"00",	-- Hex Addr	2D76	11638
x"00",	-- Hex Addr	2D77	11639
x"00",	-- Hex Addr	2D78	11640
x"00",	-- Hex Addr	2D79	11641
x"00",	-- Hex Addr	2D7A	11642
x"00",	-- Hex Addr	2D7B	11643
x"00",	-- Hex Addr	2D7C	11644
x"00",	-- Hex Addr	2D7D	11645
x"00",	-- Hex Addr	2D7E	11646
x"00",	-- Hex Addr	2D7F	11647
x"00",	-- Hex Addr	2D80	11648
x"00",	-- Hex Addr	2D81	11649
x"00",	-- Hex Addr	2D82	11650
x"00",	-- Hex Addr	2D83	11651
x"00",	-- Hex Addr	2D84	11652
x"00",	-- Hex Addr	2D85	11653
x"00",	-- Hex Addr	2D86	11654
x"00",	-- Hex Addr	2D87	11655
x"00",	-- Hex Addr	2D88	11656
x"00",	-- Hex Addr	2D89	11657
x"00",	-- Hex Addr	2D8A	11658
x"00",	-- Hex Addr	2D8B	11659
x"00",	-- Hex Addr	2D8C	11660
x"00",	-- Hex Addr	2D8D	11661
x"00",	-- Hex Addr	2D8E	11662
x"00",	-- Hex Addr	2D8F	11663
x"00",	-- Hex Addr	2D90	11664
x"00",	-- Hex Addr	2D91	11665
x"00",	-- Hex Addr	2D92	11666
x"00",	-- Hex Addr	2D93	11667
x"00",	-- Hex Addr	2D94	11668
x"00",	-- Hex Addr	2D95	11669
x"00",	-- Hex Addr	2D96	11670
x"00",	-- Hex Addr	2D97	11671
x"00",	-- Hex Addr	2D98	11672
x"00",	-- Hex Addr	2D99	11673
x"00",	-- Hex Addr	2D9A	11674
x"00",	-- Hex Addr	2D9B	11675
x"00",	-- Hex Addr	2D9C	11676
x"00",	-- Hex Addr	2D9D	11677
x"00",	-- Hex Addr	2D9E	11678
x"00",	-- Hex Addr	2D9F	11679
x"00",	-- Hex Addr	2DA0	11680
x"00",	-- Hex Addr	2DA1	11681
x"00",	-- Hex Addr	2DA2	11682
x"00",	-- Hex Addr	2DA3	11683
x"00",	-- Hex Addr	2DA4	11684
x"00",	-- Hex Addr	2DA5	11685
x"00",	-- Hex Addr	2DA6	11686
x"00",	-- Hex Addr	2DA7	11687
x"00",	-- Hex Addr	2DA8	11688
x"00",	-- Hex Addr	2DA9	11689
x"00",	-- Hex Addr	2DAA	11690
x"00",	-- Hex Addr	2DAB	11691
x"00",	-- Hex Addr	2DAC	11692
x"00",	-- Hex Addr	2DAD	11693
x"00",	-- Hex Addr	2DAE	11694
x"00",	-- Hex Addr	2DAF	11695
x"00",	-- Hex Addr	2DB0	11696
x"00",	-- Hex Addr	2DB1	11697
x"00",	-- Hex Addr	2DB2	11698
x"00",	-- Hex Addr	2DB3	11699
x"00",	-- Hex Addr	2DB4	11700
x"00",	-- Hex Addr	2DB5	11701
x"00",	-- Hex Addr	2DB6	11702
x"00",	-- Hex Addr	2DB7	11703
x"00",	-- Hex Addr	2DB8	11704
x"00",	-- Hex Addr	2DB9	11705
x"00",	-- Hex Addr	2DBA	11706
x"00",	-- Hex Addr	2DBB	11707
x"00",	-- Hex Addr	2DBC	11708
x"00",	-- Hex Addr	2DBD	11709
x"00",	-- Hex Addr	2DBE	11710
x"00",	-- Hex Addr	2DBF	11711
x"00",	-- Hex Addr	2DC0	11712
x"00",	-- Hex Addr	2DC1	11713
x"00",	-- Hex Addr	2DC2	11714
x"00",	-- Hex Addr	2DC3	11715
x"00",	-- Hex Addr	2DC4	11716
x"00",	-- Hex Addr	2DC5	11717
x"00",	-- Hex Addr	2DC6	11718
x"00",	-- Hex Addr	2DC7	11719
x"00",	-- Hex Addr	2DC8	11720
x"00",	-- Hex Addr	2DC9	11721
x"00",	-- Hex Addr	2DCA	11722
x"00",	-- Hex Addr	2DCB	11723
x"00",	-- Hex Addr	2DCC	11724
x"00",	-- Hex Addr	2DCD	11725
x"00",	-- Hex Addr	2DCE	11726
x"00",	-- Hex Addr	2DCF	11727
x"00",	-- Hex Addr	2DD0	11728
x"00",	-- Hex Addr	2DD1	11729
x"00",	-- Hex Addr	2DD2	11730
x"00",	-- Hex Addr	2DD3	11731
x"00",	-- Hex Addr	2DD4	11732
x"00",	-- Hex Addr	2DD5	11733
x"00",	-- Hex Addr	2DD6	11734
x"00",	-- Hex Addr	2DD7	11735
x"00",	-- Hex Addr	2DD8	11736
x"00",	-- Hex Addr	2DD9	11737
x"00",	-- Hex Addr	2DDA	11738
x"00",	-- Hex Addr	2DDB	11739
x"00",	-- Hex Addr	2DDC	11740
x"00",	-- Hex Addr	2DDD	11741
x"00",	-- Hex Addr	2DDE	11742
x"00",	-- Hex Addr	2DDF	11743
x"00",	-- Hex Addr	2DE0	11744
x"00",	-- Hex Addr	2DE1	11745
x"00",	-- Hex Addr	2DE2	11746
x"00",	-- Hex Addr	2DE3	11747
x"00",	-- Hex Addr	2DE4	11748
x"00",	-- Hex Addr	2DE5	11749
x"00",	-- Hex Addr	2DE6	11750
x"00",	-- Hex Addr	2DE7	11751
x"00",	-- Hex Addr	2DE8	11752
x"00",	-- Hex Addr	2DE9	11753
x"00",	-- Hex Addr	2DEA	11754
x"00",	-- Hex Addr	2DEB	11755
x"00",	-- Hex Addr	2DEC	11756
x"00",	-- Hex Addr	2DED	11757
x"00",	-- Hex Addr	2DEE	11758
x"00",	-- Hex Addr	2DEF	11759
x"00",	-- Hex Addr	2DF0	11760
x"00",	-- Hex Addr	2DF1	11761
x"00",	-- Hex Addr	2DF2	11762
x"00",	-- Hex Addr	2DF3	11763
x"00",	-- Hex Addr	2DF4	11764
x"00",	-- Hex Addr	2DF5	11765
x"00",	-- Hex Addr	2DF6	11766
x"00",	-- Hex Addr	2DF7	11767
x"00",	-- Hex Addr	2DF8	11768
x"00",	-- Hex Addr	2DF9	11769
x"00",	-- Hex Addr	2DFA	11770
x"00",	-- Hex Addr	2DFB	11771
x"00",	-- Hex Addr	2DFC	11772
x"00",	-- Hex Addr	2DFD	11773
x"00",	-- Hex Addr	2DFE	11774
x"00",	-- Hex Addr	2DFF	11775
x"00",	-- Hex Addr	2E00	11776
x"00",	-- Hex Addr	2E01	11777
x"00",	-- Hex Addr	2E02	11778
x"00",	-- Hex Addr	2E03	11779
x"00",	-- Hex Addr	2E04	11780
x"00",	-- Hex Addr	2E05	11781
x"00",	-- Hex Addr	2E06	11782
x"00",	-- Hex Addr	2E07	11783
x"00",	-- Hex Addr	2E08	11784
x"00",	-- Hex Addr	2E09	11785
x"00",	-- Hex Addr	2E0A	11786
x"00",	-- Hex Addr	2E0B	11787
x"00",	-- Hex Addr	2E0C	11788
x"00",	-- Hex Addr	2E0D	11789
x"00",	-- Hex Addr	2E0E	11790
x"00",	-- Hex Addr	2E0F	11791
x"00",	-- Hex Addr	2E10	11792
x"00",	-- Hex Addr	2E11	11793
x"00",	-- Hex Addr	2E12	11794
x"00",	-- Hex Addr	2E13	11795
x"00",	-- Hex Addr	2E14	11796
x"00",	-- Hex Addr	2E15	11797
x"00",	-- Hex Addr	2E16	11798
x"00",	-- Hex Addr	2E17	11799
x"00",	-- Hex Addr	2E18	11800
x"00",	-- Hex Addr	2E19	11801
x"00",	-- Hex Addr	2E1A	11802
x"00",	-- Hex Addr	2E1B	11803
x"00",	-- Hex Addr	2E1C	11804
x"00",	-- Hex Addr	2E1D	11805
x"00",	-- Hex Addr	2E1E	11806
x"00",	-- Hex Addr	2E1F	11807
x"00",	-- Hex Addr	2E20	11808
x"00",	-- Hex Addr	2E21	11809
x"00",	-- Hex Addr	2E22	11810
x"00",	-- Hex Addr	2E23	11811
x"00",	-- Hex Addr	2E24	11812
x"00",	-- Hex Addr	2E25	11813
x"00",	-- Hex Addr	2E26	11814
x"00",	-- Hex Addr	2E27	11815
x"00",	-- Hex Addr	2E28	11816
x"00",	-- Hex Addr	2E29	11817
x"00",	-- Hex Addr	2E2A	11818
x"00",	-- Hex Addr	2E2B	11819
x"00",	-- Hex Addr	2E2C	11820
x"00",	-- Hex Addr	2E2D	11821
x"00",	-- Hex Addr	2E2E	11822
x"00",	-- Hex Addr	2E2F	11823
x"00",	-- Hex Addr	2E30	11824
x"00",	-- Hex Addr	2E31	11825
x"00",	-- Hex Addr	2E32	11826
x"00",	-- Hex Addr	2E33	11827
x"00",	-- Hex Addr	2E34	11828
x"00",	-- Hex Addr	2E35	11829
x"00",	-- Hex Addr	2E36	11830
x"00",	-- Hex Addr	2E37	11831
x"00",	-- Hex Addr	2E38	11832
x"00",	-- Hex Addr	2E39	11833
x"00",	-- Hex Addr	2E3A	11834
x"00",	-- Hex Addr	2E3B	11835
x"00",	-- Hex Addr	2E3C	11836
x"00",	-- Hex Addr	2E3D	11837
x"00",	-- Hex Addr	2E3E	11838
x"00",	-- Hex Addr	2E3F	11839
x"00",	-- Hex Addr	2E40	11840
x"00",	-- Hex Addr	2E41	11841
x"00",	-- Hex Addr	2E42	11842
x"00",	-- Hex Addr	2E43	11843
x"00",	-- Hex Addr	2E44	11844
x"00",	-- Hex Addr	2E45	11845
x"00",	-- Hex Addr	2E46	11846
x"00",	-- Hex Addr	2E47	11847
x"00",	-- Hex Addr	2E48	11848
x"00",	-- Hex Addr	2E49	11849
x"00",	-- Hex Addr	2E4A	11850
x"00",	-- Hex Addr	2E4B	11851
x"00",	-- Hex Addr	2E4C	11852
x"00",	-- Hex Addr	2E4D	11853
x"00",	-- Hex Addr	2E4E	11854
x"00",	-- Hex Addr	2E4F	11855
x"00",	-- Hex Addr	2E50	11856
x"00",	-- Hex Addr	2E51	11857
x"00",	-- Hex Addr	2E52	11858
x"00",	-- Hex Addr	2E53	11859
x"00",	-- Hex Addr	2E54	11860
x"00",	-- Hex Addr	2E55	11861
x"00",	-- Hex Addr	2E56	11862
x"00",	-- Hex Addr	2E57	11863
x"00",	-- Hex Addr	2E58	11864
x"00",	-- Hex Addr	2E59	11865
x"00",	-- Hex Addr	2E5A	11866
x"00",	-- Hex Addr	2E5B	11867
x"00",	-- Hex Addr	2E5C	11868
x"00",	-- Hex Addr	2E5D	11869
x"00",	-- Hex Addr	2E5E	11870
x"00",	-- Hex Addr	2E5F	11871
x"00",	-- Hex Addr	2E60	11872
x"00",	-- Hex Addr	2E61	11873
x"00",	-- Hex Addr	2E62	11874
x"00",	-- Hex Addr	2E63	11875
x"00",	-- Hex Addr	2E64	11876
x"00",	-- Hex Addr	2E65	11877
x"00",	-- Hex Addr	2E66	11878
x"00",	-- Hex Addr	2E67	11879
x"00",	-- Hex Addr	2E68	11880
x"00",	-- Hex Addr	2E69	11881
x"00",	-- Hex Addr	2E6A	11882
x"00",	-- Hex Addr	2E6B	11883
x"00",	-- Hex Addr	2E6C	11884
x"00",	-- Hex Addr	2E6D	11885
x"00",	-- Hex Addr	2E6E	11886
x"00",	-- Hex Addr	2E6F	11887
x"00",	-- Hex Addr	2E70	11888
x"00",	-- Hex Addr	2E71	11889
x"00",	-- Hex Addr	2E72	11890
x"00",	-- Hex Addr	2E73	11891
x"00",	-- Hex Addr	2E74	11892
x"00",	-- Hex Addr	2E75	11893
x"00",	-- Hex Addr	2E76	11894
x"00",	-- Hex Addr	2E77	11895
x"00",	-- Hex Addr	2E78	11896
x"00",	-- Hex Addr	2E79	11897
x"00",	-- Hex Addr	2E7A	11898
x"00",	-- Hex Addr	2E7B	11899
x"00",	-- Hex Addr	2E7C	11900
x"00",	-- Hex Addr	2E7D	11901
x"00",	-- Hex Addr	2E7E	11902
x"00",	-- Hex Addr	2E7F	11903
x"00",	-- Hex Addr	2E80	11904
x"00",	-- Hex Addr	2E81	11905
x"00",	-- Hex Addr	2E82	11906
x"00",	-- Hex Addr	2E83	11907
x"00",	-- Hex Addr	2E84	11908
x"00",	-- Hex Addr	2E85	11909
x"00",	-- Hex Addr	2E86	11910
x"00",	-- Hex Addr	2E87	11911
x"00",	-- Hex Addr	2E88	11912
x"00",	-- Hex Addr	2E89	11913
x"00",	-- Hex Addr	2E8A	11914
x"00",	-- Hex Addr	2E8B	11915
x"00",	-- Hex Addr	2E8C	11916
x"00",	-- Hex Addr	2E8D	11917
x"00",	-- Hex Addr	2E8E	11918
x"00",	-- Hex Addr	2E8F	11919
x"00",	-- Hex Addr	2E90	11920
x"00",	-- Hex Addr	2E91	11921
x"00",	-- Hex Addr	2E92	11922
x"00",	-- Hex Addr	2E93	11923
x"00",	-- Hex Addr	2E94	11924
x"00",	-- Hex Addr	2E95	11925
x"00",	-- Hex Addr	2E96	11926
x"00",	-- Hex Addr	2E97	11927
x"00",	-- Hex Addr	2E98	11928
x"00",	-- Hex Addr	2E99	11929
x"00",	-- Hex Addr	2E9A	11930
x"00",	-- Hex Addr	2E9B	11931
x"00",	-- Hex Addr	2E9C	11932
x"00",	-- Hex Addr	2E9D	11933
x"00",	-- Hex Addr	2E9E	11934
x"00",	-- Hex Addr	2E9F	11935
x"00",	-- Hex Addr	2EA0	11936
x"00",	-- Hex Addr	2EA1	11937
x"00",	-- Hex Addr	2EA2	11938
x"00",	-- Hex Addr	2EA3	11939
x"00",	-- Hex Addr	2EA4	11940
x"00",	-- Hex Addr	2EA5	11941
x"00",	-- Hex Addr	2EA6	11942
x"00",	-- Hex Addr	2EA7	11943
x"00",	-- Hex Addr	2EA8	11944
x"00",	-- Hex Addr	2EA9	11945
x"00",	-- Hex Addr	2EAA	11946
x"00",	-- Hex Addr	2EAB	11947
x"00",	-- Hex Addr	2EAC	11948
x"00",	-- Hex Addr	2EAD	11949
x"00",	-- Hex Addr	2EAE	11950
x"00",	-- Hex Addr	2EAF	11951
x"00",	-- Hex Addr	2EB0	11952
x"00",	-- Hex Addr	2EB1	11953
x"00",	-- Hex Addr	2EB2	11954
x"00",	-- Hex Addr	2EB3	11955
x"00",	-- Hex Addr	2EB4	11956
x"00",	-- Hex Addr	2EB5	11957
x"00",	-- Hex Addr	2EB6	11958
x"00",	-- Hex Addr	2EB7	11959
x"00",	-- Hex Addr	2EB8	11960
x"00",	-- Hex Addr	2EB9	11961
x"00",	-- Hex Addr	2EBA	11962
x"00",	-- Hex Addr	2EBB	11963
x"00",	-- Hex Addr	2EBC	11964
x"00",	-- Hex Addr	2EBD	11965
x"00",	-- Hex Addr	2EBE	11966
x"00",	-- Hex Addr	2EBF	11967
x"00",	-- Hex Addr	2EC0	11968
x"00",	-- Hex Addr	2EC1	11969
x"00",	-- Hex Addr	2EC2	11970
x"00",	-- Hex Addr	2EC3	11971
x"00",	-- Hex Addr	2EC4	11972
x"00",	-- Hex Addr	2EC5	11973
x"00",	-- Hex Addr	2EC6	11974
x"00",	-- Hex Addr	2EC7	11975
x"00",	-- Hex Addr	2EC8	11976
x"00",	-- Hex Addr	2EC9	11977
x"00",	-- Hex Addr	2ECA	11978
x"00",	-- Hex Addr	2ECB	11979
x"00",	-- Hex Addr	2ECC	11980
x"00",	-- Hex Addr	2ECD	11981
x"00",	-- Hex Addr	2ECE	11982
x"00",	-- Hex Addr	2ECF	11983
x"00",	-- Hex Addr	2ED0	11984
x"00",	-- Hex Addr	2ED1	11985
x"00",	-- Hex Addr	2ED2	11986
x"00",	-- Hex Addr	2ED3	11987
x"00",	-- Hex Addr	2ED4	11988
x"00",	-- Hex Addr	2ED5	11989
x"00",	-- Hex Addr	2ED6	11990
x"00",	-- Hex Addr	2ED7	11991
x"00",	-- Hex Addr	2ED8	11992
x"00",	-- Hex Addr	2ED9	11993
x"00",	-- Hex Addr	2EDA	11994
x"00",	-- Hex Addr	2EDB	11995
x"00",	-- Hex Addr	2EDC	11996
x"00",	-- Hex Addr	2EDD	11997
x"00",	-- Hex Addr	2EDE	11998
x"00",	-- Hex Addr	2EDF	11999
x"00",	-- Hex Addr	2EE0	12000
x"00",	-- Hex Addr	2EE1	12001
x"00",	-- Hex Addr	2EE2	12002
x"00",	-- Hex Addr	2EE3	12003
x"00",	-- Hex Addr	2EE4	12004
x"00",	-- Hex Addr	2EE5	12005
x"00",	-- Hex Addr	2EE6	12006
x"00",	-- Hex Addr	2EE7	12007
x"00",	-- Hex Addr	2EE8	12008
x"00",	-- Hex Addr	2EE9	12009
x"00",	-- Hex Addr	2EEA	12010
x"00",	-- Hex Addr	2EEB	12011
x"00",	-- Hex Addr	2EEC	12012
x"00",	-- Hex Addr	2EED	12013
x"00",	-- Hex Addr	2EEE	12014
x"00",	-- Hex Addr	2EEF	12015
x"00",	-- Hex Addr	2EF0	12016
x"00",	-- Hex Addr	2EF1	12017
x"00",	-- Hex Addr	2EF2	12018
x"00",	-- Hex Addr	2EF3	12019
x"00",	-- Hex Addr	2EF4	12020
x"00",	-- Hex Addr	2EF5	12021
x"00",	-- Hex Addr	2EF6	12022
x"00",	-- Hex Addr	2EF7	12023
x"00",	-- Hex Addr	2EF8	12024
x"00",	-- Hex Addr	2EF9	12025
x"00",	-- Hex Addr	2EFA	12026
x"00",	-- Hex Addr	2EFB	12027
x"00",	-- Hex Addr	2EFC	12028
x"00",	-- Hex Addr	2EFD	12029
x"00",	-- Hex Addr	2EFE	12030
x"00",	-- Hex Addr	2EFF	12031
x"00",	-- Hex Addr	2F00	12032
x"00",	-- Hex Addr	2F01	12033
x"00",	-- Hex Addr	2F02	12034
x"00",	-- Hex Addr	2F03	12035
x"00",	-- Hex Addr	2F04	12036
x"00",	-- Hex Addr	2F05	12037
x"00",	-- Hex Addr	2F06	12038
x"00",	-- Hex Addr	2F07	12039
x"00",	-- Hex Addr	2F08	12040
x"00",	-- Hex Addr	2F09	12041
x"00",	-- Hex Addr	2F0A	12042
x"00",	-- Hex Addr	2F0B	12043
x"00",	-- Hex Addr	2F0C	12044
x"00",	-- Hex Addr	2F0D	12045
x"00",	-- Hex Addr	2F0E	12046
x"00",	-- Hex Addr	2F0F	12047
x"00",	-- Hex Addr	2F10	12048
x"00",	-- Hex Addr	2F11	12049
x"00",	-- Hex Addr	2F12	12050
x"00",	-- Hex Addr	2F13	12051
x"00",	-- Hex Addr	2F14	12052
x"00",	-- Hex Addr	2F15	12053
x"00",	-- Hex Addr	2F16	12054
x"00",	-- Hex Addr	2F17	12055
x"00",	-- Hex Addr	2F18	12056
x"00",	-- Hex Addr	2F19	12057
x"00",	-- Hex Addr	2F1A	12058
x"00",	-- Hex Addr	2F1B	12059
x"00",	-- Hex Addr	2F1C	12060
x"00",	-- Hex Addr	2F1D	12061
x"00",	-- Hex Addr	2F1E	12062
x"00",	-- Hex Addr	2F1F	12063
x"00",	-- Hex Addr	2F20	12064
x"00",	-- Hex Addr	2F21	12065
x"00",	-- Hex Addr	2F22	12066
x"00",	-- Hex Addr	2F23	12067
x"00",	-- Hex Addr	2F24	12068
x"00",	-- Hex Addr	2F25	12069
x"00",	-- Hex Addr	2F26	12070
x"00",	-- Hex Addr	2F27	12071
x"00",	-- Hex Addr	2F28	12072
x"00",	-- Hex Addr	2F29	12073
x"00",	-- Hex Addr	2F2A	12074
x"00",	-- Hex Addr	2F2B	12075
x"00",	-- Hex Addr	2F2C	12076
x"00",	-- Hex Addr	2F2D	12077
x"00",	-- Hex Addr	2F2E	12078
x"00",	-- Hex Addr	2F2F	12079
x"00",	-- Hex Addr	2F30	12080
x"00",	-- Hex Addr	2F31	12081
x"00",	-- Hex Addr	2F32	12082
x"00",	-- Hex Addr	2F33	12083
x"00",	-- Hex Addr	2F34	12084
x"00",	-- Hex Addr	2F35	12085
x"00",	-- Hex Addr	2F36	12086
x"00",	-- Hex Addr	2F37	12087
x"00",	-- Hex Addr	2F38	12088
x"00",	-- Hex Addr	2F39	12089
x"00",	-- Hex Addr	2F3A	12090
x"00",	-- Hex Addr	2F3B	12091
x"00",	-- Hex Addr	2F3C	12092
x"00",	-- Hex Addr	2F3D	12093
x"00",	-- Hex Addr	2F3E	12094
x"00",	-- Hex Addr	2F3F	12095
x"00",	-- Hex Addr	2F40	12096
x"00",	-- Hex Addr	2F41	12097
x"00",	-- Hex Addr	2F42	12098
x"00",	-- Hex Addr	2F43	12099
x"00",	-- Hex Addr	2F44	12100
x"00",	-- Hex Addr	2F45	12101
x"00",	-- Hex Addr	2F46	12102
x"00",	-- Hex Addr	2F47	12103
x"00",	-- Hex Addr	2F48	12104
x"00",	-- Hex Addr	2F49	12105
x"00",	-- Hex Addr	2F4A	12106
x"00",	-- Hex Addr	2F4B	12107
x"00",	-- Hex Addr	2F4C	12108
x"00",	-- Hex Addr	2F4D	12109
x"00",	-- Hex Addr	2F4E	12110
x"00",	-- Hex Addr	2F4F	12111
x"00",	-- Hex Addr	2F50	12112
x"00",	-- Hex Addr	2F51	12113
x"00",	-- Hex Addr	2F52	12114
x"00",	-- Hex Addr	2F53	12115
x"00",	-- Hex Addr	2F54	12116
x"00",	-- Hex Addr	2F55	12117
x"00",	-- Hex Addr	2F56	12118
x"00",	-- Hex Addr	2F57	12119
x"00",	-- Hex Addr	2F58	12120
x"00",	-- Hex Addr	2F59	12121
x"00",	-- Hex Addr	2F5A	12122
x"00",	-- Hex Addr	2F5B	12123
x"00",	-- Hex Addr	2F5C	12124
x"00",	-- Hex Addr	2F5D	12125
x"00",	-- Hex Addr	2F5E	12126
x"00",	-- Hex Addr	2F5F	12127
x"00",	-- Hex Addr	2F60	12128
x"00",	-- Hex Addr	2F61	12129
x"00",	-- Hex Addr	2F62	12130
x"00",	-- Hex Addr	2F63	12131
x"00",	-- Hex Addr	2F64	12132
x"00",	-- Hex Addr	2F65	12133
x"00",	-- Hex Addr	2F66	12134
x"00",	-- Hex Addr	2F67	12135
x"00",	-- Hex Addr	2F68	12136
x"00",	-- Hex Addr	2F69	12137
x"00",	-- Hex Addr	2F6A	12138
x"00",	-- Hex Addr	2F6B	12139
x"00",	-- Hex Addr	2F6C	12140
x"00",	-- Hex Addr	2F6D	12141
x"00",	-- Hex Addr	2F6E	12142
x"00",	-- Hex Addr	2F6F	12143
x"00",	-- Hex Addr	2F70	12144
x"00",	-- Hex Addr	2F71	12145
x"00",	-- Hex Addr	2F72	12146
x"00",	-- Hex Addr	2F73	12147
x"00",	-- Hex Addr	2F74	12148
x"00",	-- Hex Addr	2F75	12149
x"00",	-- Hex Addr	2F76	12150
x"00",	-- Hex Addr	2F77	12151
x"00",	-- Hex Addr	2F78	12152
x"00",	-- Hex Addr	2F79	12153
x"00",	-- Hex Addr	2F7A	12154
x"00",	-- Hex Addr	2F7B	12155
x"00",	-- Hex Addr	2F7C	12156
x"00",	-- Hex Addr	2F7D	12157
x"00",	-- Hex Addr	2F7E	12158
x"00",	-- Hex Addr	2F7F	12159
x"00",	-- Hex Addr	2F80	12160
x"00",	-- Hex Addr	2F81	12161
x"00",	-- Hex Addr	2F82	12162
x"00",	-- Hex Addr	2F83	12163
x"00",	-- Hex Addr	2F84	12164
x"00",	-- Hex Addr	2F85	12165
x"00",	-- Hex Addr	2F86	12166
x"00",	-- Hex Addr	2F87	12167
x"00",	-- Hex Addr	2F88	12168
x"00",	-- Hex Addr	2F89	12169
x"00",	-- Hex Addr	2F8A	12170
x"00",	-- Hex Addr	2F8B	12171
x"00",	-- Hex Addr	2F8C	12172
x"00",	-- Hex Addr	2F8D	12173
x"00",	-- Hex Addr	2F8E	12174
x"00",	-- Hex Addr	2F8F	12175
x"00",	-- Hex Addr	2F90	12176
x"00",	-- Hex Addr	2F91	12177
x"00",	-- Hex Addr	2F92	12178
x"00",	-- Hex Addr	2F93	12179
x"00",	-- Hex Addr	2F94	12180
x"00",	-- Hex Addr	2F95	12181
x"00",	-- Hex Addr	2F96	12182
x"00",	-- Hex Addr	2F97	12183
x"00",	-- Hex Addr	2F98	12184
x"00",	-- Hex Addr	2F99	12185
x"00",	-- Hex Addr	2F9A	12186
x"00",	-- Hex Addr	2F9B	12187
x"00",	-- Hex Addr	2F9C	12188
x"00",	-- Hex Addr	2F9D	12189
x"00",	-- Hex Addr	2F9E	12190
x"00",	-- Hex Addr	2F9F	12191
x"00",	-- Hex Addr	2FA0	12192
x"00",	-- Hex Addr	2FA1	12193
x"00",	-- Hex Addr	2FA2	12194
x"00",	-- Hex Addr	2FA3	12195
x"00",	-- Hex Addr	2FA4	12196
x"00",	-- Hex Addr	2FA5	12197
x"00",	-- Hex Addr	2FA6	12198
x"00",	-- Hex Addr	2FA7	12199
x"00",	-- Hex Addr	2FA8	12200
x"00",	-- Hex Addr	2FA9	12201
x"00",	-- Hex Addr	2FAA	12202
x"00",	-- Hex Addr	2FAB	12203
x"00",	-- Hex Addr	2FAC	12204
x"00",	-- Hex Addr	2FAD	12205
x"00",	-- Hex Addr	2FAE	12206
x"00",	-- Hex Addr	2FAF	12207
x"00",	-- Hex Addr	2FB0	12208
x"00",	-- Hex Addr	2FB1	12209
x"00",	-- Hex Addr	2FB2	12210
x"00",	-- Hex Addr	2FB3	12211
x"00",	-- Hex Addr	2FB4	12212
x"00",	-- Hex Addr	2FB5	12213
x"00",	-- Hex Addr	2FB6	12214
x"00",	-- Hex Addr	2FB7	12215
x"00",	-- Hex Addr	2FB8	12216
x"00",	-- Hex Addr	2FB9	12217
x"00",	-- Hex Addr	2FBA	12218
x"00",	-- Hex Addr	2FBB	12219
x"00",	-- Hex Addr	2FBC	12220
x"00",	-- Hex Addr	2FBD	12221
x"00",	-- Hex Addr	2FBE	12222
x"00",	-- Hex Addr	2FBF	12223
x"00",	-- Hex Addr	2FC0	12224
x"00",	-- Hex Addr	2FC1	12225
x"00",	-- Hex Addr	2FC2	12226
x"00",	-- Hex Addr	2FC3	12227
x"00",	-- Hex Addr	2FC4	12228
x"00",	-- Hex Addr	2FC5	12229
x"00",	-- Hex Addr	2FC6	12230
x"00",	-- Hex Addr	2FC7	12231
x"00",	-- Hex Addr	2FC8	12232
x"00",	-- Hex Addr	2FC9	12233
x"00",	-- Hex Addr	2FCA	12234
x"00",	-- Hex Addr	2FCB	12235
x"00",	-- Hex Addr	2FCC	12236
x"00",	-- Hex Addr	2FCD	12237
x"00",	-- Hex Addr	2FCE	12238
x"00",	-- Hex Addr	2FCF	12239
x"00",	-- Hex Addr	2FD0	12240
x"00",	-- Hex Addr	2FD1	12241
x"00",	-- Hex Addr	2FD2	12242
x"00",	-- Hex Addr	2FD3	12243
x"00",	-- Hex Addr	2FD4	12244
x"00",	-- Hex Addr	2FD5	12245
x"00",	-- Hex Addr	2FD6	12246
x"00",	-- Hex Addr	2FD7	12247
x"00",	-- Hex Addr	2FD8	12248
x"00",	-- Hex Addr	2FD9	12249
x"00",	-- Hex Addr	2FDA	12250
x"00",	-- Hex Addr	2FDB	12251
x"00",	-- Hex Addr	2FDC	12252
x"00",	-- Hex Addr	2FDD	12253
x"00",	-- Hex Addr	2FDE	12254
x"00",	-- Hex Addr	2FDF	12255
x"00",	-- Hex Addr	2FE0	12256
x"00",	-- Hex Addr	2FE1	12257
x"00",	-- Hex Addr	2FE2	12258
x"00",	-- Hex Addr	2FE3	12259
x"00",	-- Hex Addr	2FE4	12260
x"00",	-- Hex Addr	2FE5	12261
x"00",	-- Hex Addr	2FE6	12262
x"00",	-- Hex Addr	2FE7	12263
x"00",	-- Hex Addr	2FE8	12264
x"00",	-- Hex Addr	2FE9	12265
x"00",	-- Hex Addr	2FEA	12266
x"00",	-- Hex Addr	2FEB	12267
x"00",	-- Hex Addr	2FEC	12268
x"00",	-- Hex Addr	2FED	12269
x"00",	-- Hex Addr	2FEE	12270
x"00",	-- Hex Addr	2FEF	12271
x"00",	-- Hex Addr	2FF0	12272
x"00",	-- Hex Addr	2FF1	12273
x"00",	-- Hex Addr	2FF2	12274
x"00",	-- Hex Addr	2FF3	12275
x"00",	-- Hex Addr	2FF4	12276
x"00",	-- Hex Addr	2FF5	12277
x"00",	-- Hex Addr	2FF6	12278
x"00",	-- Hex Addr	2FF7	12279
x"00",	-- Hex Addr	2FF8	12280
x"00",	-- Hex Addr	2FF9	12281
x"00",	-- Hex Addr	2FFA	12282
x"00",	-- Hex Addr	2FFB	12283
x"00",	-- Hex Addr	2FFC	12284
x"00",	-- Hex Addr	2FFD	12285
x"00",	-- Hex Addr	2FFE	12286
x"00",	-- Hex Addr	2FFF	12287
x"00",	-- Hex Addr	3000	12288
x"00",	-- Hex Addr	3001	12289
x"00",	-- Hex Addr	3002	12290
x"00",	-- Hex Addr	3003	12291
x"00",	-- Hex Addr	3004	12292
x"00",	-- Hex Addr	3005	12293
x"00",	-- Hex Addr	3006	12294
x"00",	-- Hex Addr	3007	12295
x"00",	-- Hex Addr	3008	12296
x"00",	-- Hex Addr	3009	12297
x"00",	-- Hex Addr	300A	12298
x"00",	-- Hex Addr	300B	12299
x"00",	-- Hex Addr	300C	12300
x"00",	-- Hex Addr	300D	12301
x"00",	-- Hex Addr	300E	12302
x"00",	-- Hex Addr	300F	12303
x"00",	-- Hex Addr	3010	12304
x"00",	-- Hex Addr	3011	12305
x"00",	-- Hex Addr	3012	12306
x"00",	-- Hex Addr	3013	12307
x"00",	-- Hex Addr	3014	12308
x"00",	-- Hex Addr	3015	12309
x"00",	-- Hex Addr	3016	12310
x"00",	-- Hex Addr	3017	12311
x"00",	-- Hex Addr	3018	12312
x"00",	-- Hex Addr	3019	12313
x"00",	-- Hex Addr	301A	12314
x"00",	-- Hex Addr	301B	12315
x"00",	-- Hex Addr	301C	12316
x"00",	-- Hex Addr	301D	12317
x"00",	-- Hex Addr	301E	12318
x"00",	-- Hex Addr	301F	12319
x"00",	-- Hex Addr	3020	12320
x"00",	-- Hex Addr	3021	12321
x"00",	-- Hex Addr	3022	12322
x"00",	-- Hex Addr	3023	12323
x"00",	-- Hex Addr	3024	12324
x"00",	-- Hex Addr	3025	12325
x"00",	-- Hex Addr	3026	12326
x"00",	-- Hex Addr	3027	12327
x"00",	-- Hex Addr	3028	12328
x"00",	-- Hex Addr	3029	12329
x"00",	-- Hex Addr	302A	12330
x"00",	-- Hex Addr	302B	12331
x"00",	-- Hex Addr	302C	12332
x"00",	-- Hex Addr	302D	12333
x"00",	-- Hex Addr	302E	12334
x"00",	-- Hex Addr	302F	12335
x"00",	-- Hex Addr	3030	12336
x"00",	-- Hex Addr	3031	12337
x"00",	-- Hex Addr	3032	12338
x"00",	-- Hex Addr	3033	12339
x"00",	-- Hex Addr	3034	12340
x"00",	-- Hex Addr	3035	12341
x"00",	-- Hex Addr	3036	12342
x"00",	-- Hex Addr	3037	12343
x"00",	-- Hex Addr	3038	12344
x"00",	-- Hex Addr	3039	12345
x"00",	-- Hex Addr	303A	12346
x"00",	-- Hex Addr	303B	12347
x"00",	-- Hex Addr	303C	12348
x"00",	-- Hex Addr	303D	12349
x"00",	-- Hex Addr	303E	12350
x"00",	-- Hex Addr	303F	12351
x"00",	-- Hex Addr	3040	12352
x"00",	-- Hex Addr	3041	12353
x"00",	-- Hex Addr	3042	12354
x"00",	-- Hex Addr	3043	12355
x"00",	-- Hex Addr	3044	12356
x"00",	-- Hex Addr	3045	12357
x"00",	-- Hex Addr	3046	12358
x"00",	-- Hex Addr	3047	12359
x"00",	-- Hex Addr	3048	12360
x"00",	-- Hex Addr	3049	12361
x"00",	-- Hex Addr	304A	12362
x"00",	-- Hex Addr	304B	12363
x"00",	-- Hex Addr	304C	12364
x"00",	-- Hex Addr	304D	12365
x"00",	-- Hex Addr	304E	12366
x"00",	-- Hex Addr	304F	12367
x"00",	-- Hex Addr	3050	12368
x"00",	-- Hex Addr	3051	12369
x"00",	-- Hex Addr	3052	12370
x"00",	-- Hex Addr	3053	12371
x"00",	-- Hex Addr	3054	12372
x"00",	-- Hex Addr	3055	12373
x"00",	-- Hex Addr	3056	12374
x"00",	-- Hex Addr	3057	12375
x"00",	-- Hex Addr	3058	12376
x"00",	-- Hex Addr	3059	12377
x"00",	-- Hex Addr	305A	12378
x"00",	-- Hex Addr	305B	12379
x"00",	-- Hex Addr	305C	12380
x"00",	-- Hex Addr	305D	12381
x"00",	-- Hex Addr	305E	12382
x"00",	-- Hex Addr	305F	12383
x"00",	-- Hex Addr	3060	12384
x"00",	-- Hex Addr	3061	12385
x"00",	-- Hex Addr	3062	12386
x"00",	-- Hex Addr	3063	12387
x"00",	-- Hex Addr	3064	12388
x"00",	-- Hex Addr	3065	12389
x"00",	-- Hex Addr	3066	12390
x"00",	-- Hex Addr	3067	12391
x"00",	-- Hex Addr	3068	12392
x"00",	-- Hex Addr	3069	12393
x"00",	-- Hex Addr	306A	12394
x"00",	-- Hex Addr	306B	12395
x"00",	-- Hex Addr	306C	12396
x"00",	-- Hex Addr	306D	12397
x"00",	-- Hex Addr	306E	12398
x"00",	-- Hex Addr	306F	12399
x"00",	-- Hex Addr	3070	12400
x"00",	-- Hex Addr	3071	12401
x"00",	-- Hex Addr	3072	12402
x"00",	-- Hex Addr	3073	12403
x"00",	-- Hex Addr	3074	12404
x"00",	-- Hex Addr	3075	12405
x"00",	-- Hex Addr	3076	12406
x"00",	-- Hex Addr	3077	12407
x"00",	-- Hex Addr	3078	12408
x"00",	-- Hex Addr	3079	12409
x"00",	-- Hex Addr	307A	12410
x"00",	-- Hex Addr	307B	12411
x"00",	-- Hex Addr	307C	12412
x"00",	-- Hex Addr	307D	12413
x"00",	-- Hex Addr	307E	12414
x"00",	-- Hex Addr	307F	12415
x"00",	-- Hex Addr	3080	12416
x"00",	-- Hex Addr	3081	12417
x"00",	-- Hex Addr	3082	12418
x"00",	-- Hex Addr	3083	12419
x"00",	-- Hex Addr	3084	12420
x"00",	-- Hex Addr	3085	12421
x"00",	-- Hex Addr	3086	12422
x"00",	-- Hex Addr	3087	12423
x"00",	-- Hex Addr	3088	12424
x"00",	-- Hex Addr	3089	12425
x"00",	-- Hex Addr	308A	12426
x"00",	-- Hex Addr	308B	12427
x"00",	-- Hex Addr	308C	12428
x"00",	-- Hex Addr	308D	12429
x"00",	-- Hex Addr	308E	12430
x"00",	-- Hex Addr	308F	12431
x"00",	-- Hex Addr	3090	12432
x"00",	-- Hex Addr	3091	12433
x"00",	-- Hex Addr	3092	12434
x"00",	-- Hex Addr	3093	12435
x"00",	-- Hex Addr	3094	12436
x"00",	-- Hex Addr	3095	12437
x"00",	-- Hex Addr	3096	12438
x"00",	-- Hex Addr	3097	12439
x"00",	-- Hex Addr	3098	12440
x"00",	-- Hex Addr	3099	12441
x"00",	-- Hex Addr	309A	12442
x"00",	-- Hex Addr	309B	12443
x"00",	-- Hex Addr	309C	12444
x"00",	-- Hex Addr	309D	12445
x"00",	-- Hex Addr	309E	12446
x"00",	-- Hex Addr	309F	12447
x"00",	-- Hex Addr	30A0	12448
x"00",	-- Hex Addr	30A1	12449
x"00",	-- Hex Addr	30A2	12450
x"00",	-- Hex Addr	30A3	12451
x"00",	-- Hex Addr	30A4	12452
x"00",	-- Hex Addr	30A5	12453
x"00",	-- Hex Addr	30A6	12454
x"00",	-- Hex Addr	30A7	12455
x"00",	-- Hex Addr	30A8	12456
x"00",	-- Hex Addr	30A9	12457
x"00",	-- Hex Addr	30AA	12458
x"00",	-- Hex Addr	30AB	12459
x"00",	-- Hex Addr	30AC	12460
x"00",	-- Hex Addr	30AD	12461
x"00",	-- Hex Addr	30AE	12462
x"00",	-- Hex Addr	30AF	12463
x"00",	-- Hex Addr	30B0	12464
x"00",	-- Hex Addr	30B1	12465
x"00",	-- Hex Addr	30B2	12466
x"00",	-- Hex Addr	30B3	12467
x"00",	-- Hex Addr	30B4	12468
x"00",	-- Hex Addr	30B5	12469
x"00",	-- Hex Addr	30B6	12470
x"00",	-- Hex Addr	30B7	12471
x"00",	-- Hex Addr	30B8	12472
x"00",	-- Hex Addr	30B9	12473
x"00",	-- Hex Addr	30BA	12474
x"00",	-- Hex Addr	30BB	12475
x"00",	-- Hex Addr	30BC	12476
x"00",	-- Hex Addr	30BD	12477
x"00",	-- Hex Addr	30BE	12478
x"00",	-- Hex Addr	30BF	12479
x"00",	-- Hex Addr	30C0	12480
x"00",	-- Hex Addr	30C1	12481
x"00",	-- Hex Addr	30C2	12482
x"00",	-- Hex Addr	30C3	12483
x"00",	-- Hex Addr	30C4	12484
x"00",	-- Hex Addr	30C5	12485
x"00",	-- Hex Addr	30C6	12486
x"00",	-- Hex Addr	30C7	12487
x"00",	-- Hex Addr	30C8	12488
x"00",	-- Hex Addr	30C9	12489
x"00",	-- Hex Addr	30CA	12490
x"00",	-- Hex Addr	30CB	12491
x"00",	-- Hex Addr	30CC	12492
x"00",	-- Hex Addr	30CD	12493
x"00",	-- Hex Addr	30CE	12494
x"00",	-- Hex Addr	30CF	12495
x"00",	-- Hex Addr	30D0	12496
x"00",	-- Hex Addr	30D1	12497
x"00",	-- Hex Addr	30D2	12498
x"00",	-- Hex Addr	30D3	12499
x"00",	-- Hex Addr	30D4	12500
x"00",	-- Hex Addr	30D5	12501
x"00",	-- Hex Addr	30D6	12502
x"00",	-- Hex Addr	30D7	12503
x"00",	-- Hex Addr	30D8	12504
x"00",	-- Hex Addr	30D9	12505
x"00",	-- Hex Addr	30DA	12506
x"00",	-- Hex Addr	30DB	12507
x"00",	-- Hex Addr	30DC	12508
x"00",	-- Hex Addr	30DD	12509
x"00",	-- Hex Addr	30DE	12510
x"00",	-- Hex Addr	30DF	12511
x"00",	-- Hex Addr	30E0	12512
x"00",	-- Hex Addr	30E1	12513
x"00",	-- Hex Addr	30E2	12514
x"00",	-- Hex Addr	30E3	12515
x"00",	-- Hex Addr	30E4	12516
x"00",	-- Hex Addr	30E5	12517
x"00",	-- Hex Addr	30E6	12518
x"00",	-- Hex Addr	30E7	12519
x"00",	-- Hex Addr	30E8	12520
x"00",	-- Hex Addr	30E9	12521
x"00",	-- Hex Addr	30EA	12522
x"00",	-- Hex Addr	30EB	12523
x"00",	-- Hex Addr	30EC	12524
x"00",	-- Hex Addr	30ED	12525
x"00",	-- Hex Addr	30EE	12526
x"00",	-- Hex Addr	30EF	12527
x"00",	-- Hex Addr	30F0	12528
x"00",	-- Hex Addr	30F1	12529
x"00",	-- Hex Addr	30F2	12530
x"00",	-- Hex Addr	30F3	12531
x"00",	-- Hex Addr	30F4	12532
x"00",	-- Hex Addr	30F5	12533
x"00",	-- Hex Addr	30F6	12534
x"00",	-- Hex Addr	30F7	12535
x"00",	-- Hex Addr	30F8	12536
x"00",	-- Hex Addr	30F9	12537
x"00",	-- Hex Addr	30FA	12538
x"00",	-- Hex Addr	30FB	12539
x"00",	-- Hex Addr	30FC	12540
x"00",	-- Hex Addr	30FD	12541
x"00",	-- Hex Addr	30FE	12542
x"00",	-- Hex Addr	30FF	12543
x"00",	-- Hex Addr	3100	12544
x"00",	-- Hex Addr	3101	12545
x"00",	-- Hex Addr	3102	12546
x"00",	-- Hex Addr	3103	12547
x"00",	-- Hex Addr	3104	12548
x"00",	-- Hex Addr	3105	12549
x"00",	-- Hex Addr	3106	12550
x"00",	-- Hex Addr	3107	12551
x"00",	-- Hex Addr	3108	12552
x"00",	-- Hex Addr	3109	12553
x"00",	-- Hex Addr	310A	12554
x"00",	-- Hex Addr	310B	12555
x"00",	-- Hex Addr	310C	12556
x"00",	-- Hex Addr	310D	12557
x"00",	-- Hex Addr	310E	12558
x"00",	-- Hex Addr	310F	12559
x"00",	-- Hex Addr	3110	12560
x"00",	-- Hex Addr	3111	12561
x"00",	-- Hex Addr	3112	12562
x"00",	-- Hex Addr	3113	12563
x"00",	-- Hex Addr	3114	12564
x"00",	-- Hex Addr	3115	12565
x"00",	-- Hex Addr	3116	12566
x"00",	-- Hex Addr	3117	12567
x"00",	-- Hex Addr	3118	12568
x"00",	-- Hex Addr	3119	12569
x"00",	-- Hex Addr	311A	12570
x"00",	-- Hex Addr	311B	12571
x"00",	-- Hex Addr	311C	12572
x"00",	-- Hex Addr	311D	12573
x"00",	-- Hex Addr	311E	12574
x"00",	-- Hex Addr	311F	12575
x"00",	-- Hex Addr	3120	12576
x"00",	-- Hex Addr	3121	12577
x"00",	-- Hex Addr	3122	12578
x"00",	-- Hex Addr	3123	12579
x"00",	-- Hex Addr	3124	12580
x"00",	-- Hex Addr	3125	12581
x"00",	-- Hex Addr	3126	12582
x"00",	-- Hex Addr	3127	12583
x"00",	-- Hex Addr	3128	12584
x"00",	-- Hex Addr	3129	12585
x"00",	-- Hex Addr	312A	12586
x"00",	-- Hex Addr	312B	12587
x"00",	-- Hex Addr	312C	12588
x"00",	-- Hex Addr	312D	12589
x"00",	-- Hex Addr	312E	12590
x"00",	-- Hex Addr	312F	12591
x"00",	-- Hex Addr	3130	12592
x"00",	-- Hex Addr	3131	12593
x"00",	-- Hex Addr	3132	12594
x"00",	-- Hex Addr	3133	12595
x"00",	-- Hex Addr	3134	12596
x"00",	-- Hex Addr	3135	12597
x"00",	-- Hex Addr	3136	12598
x"00",	-- Hex Addr	3137	12599
x"00",	-- Hex Addr	3138	12600
x"00",	-- Hex Addr	3139	12601
x"00",	-- Hex Addr	313A	12602
x"00",	-- Hex Addr	313B	12603
x"00",	-- Hex Addr	313C	12604
x"00",	-- Hex Addr	313D	12605
x"00",	-- Hex Addr	313E	12606
x"00",	-- Hex Addr	313F	12607
x"00",	-- Hex Addr	3140	12608
x"00",	-- Hex Addr	3141	12609
x"00",	-- Hex Addr	3142	12610
x"00",	-- Hex Addr	3143	12611
x"00",	-- Hex Addr	3144	12612
x"00",	-- Hex Addr	3145	12613
x"00",	-- Hex Addr	3146	12614
x"00",	-- Hex Addr	3147	12615
x"00",	-- Hex Addr	3148	12616
x"00",	-- Hex Addr	3149	12617
x"00",	-- Hex Addr	314A	12618
x"00",	-- Hex Addr	314B	12619
x"00",	-- Hex Addr	314C	12620
x"00",	-- Hex Addr	314D	12621
x"00",	-- Hex Addr	314E	12622
x"00",	-- Hex Addr	314F	12623
x"00",	-- Hex Addr	3150	12624
x"00",	-- Hex Addr	3151	12625
x"00",	-- Hex Addr	3152	12626
x"00",	-- Hex Addr	3153	12627
x"00",	-- Hex Addr	3154	12628
x"00",	-- Hex Addr	3155	12629
x"00",	-- Hex Addr	3156	12630
x"00",	-- Hex Addr	3157	12631
x"00",	-- Hex Addr	3158	12632
x"00",	-- Hex Addr	3159	12633
x"00",	-- Hex Addr	315A	12634
x"00",	-- Hex Addr	315B	12635
x"00",	-- Hex Addr	315C	12636
x"00",	-- Hex Addr	315D	12637
x"00",	-- Hex Addr	315E	12638
x"00",	-- Hex Addr	315F	12639
x"00",	-- Hex Addr	3160	12640
x"00",	-- Hex Addr	3161	12641
x"00",	-- Hex Addr	3162	12642
x"00",	-- Hex Addr	3163	12643
x"00",	-- Hex Addr	3164	12644
x"00",	-- Hex Addr	3165	12645
x"00",	-- Hex Addr	3166	12646
x"00",	-- Hex Addr	3167	12647
x"00",	-- Hex Addr	3168	12648
x"00",	-- Hex Addr	3169	12649
x"00",	-- Hex Addr	316A	12650
x"00",	-- Hex Addr	316B	12651
x"00",	-- Hex Addr	316C	12652
x"00",	-- Hex Addr	316D	12653
x"00",	-- Hex Addr	316E	12654
x"00",	-- Hex Addr	316F	12655
x"00",	-- Hex Addr	3170	12656
x"00",	-- Hex Addr	3171	12657
x"00",	-- Hex Addr	3172	12658
x"00",	-- Hex Addr	3173	12659
x"00",	-- Hex Addr	3174	12660
x"00",	-- Hex Addr	3175	12661
x"00",	-- Hex Addr	3176	12662
x"00",	-- Hex Addr	3177	12663
x"00",	-- Hex Addr	3178	12664
x"00",	-- Hex Addr	3179	12665
x"00",	-- Hex Addr	317A	12666
x"00",	-- Hex Addr	317B	12667
x"00",	-- Hex Addr	317C	12668
x"00",	-- Hex Addr	317D	12669
x"00",	-- Hex Addr	317E	12670
x"00",	-- Hex Addr	317F	12671
x"00",	-- Hex Addr	3180	12672
x"00",	-- Hex Addr	3181	12673
x"00",	-- Hex Addr	3182	12674
x"00",	-- Hex Addr	3183	12675
x"00",	-- Hex Addr	3184	12676
x"00",	-- Hex Addr	3185	12677
x"00",	-- Hex Addr	3186	12678
x"00",	-- Hex Addr	3187	12679
x"00",	-- Hex Addr	3188	12680
x"00",	-- Hex Addr	3189	12681
x"00",	-- Hex Addr	318A	12682
x"00",	-- Hex Addr	318B	12683
x"00",	-- Hex Addr	318C	12684
x"00",	-- Hex Addr	318D	12685
x"00",	-- Hex Addr	318E	12686
x"00",	-- Hex Addr	318F	12687
x"00",	-- Hex Addr	3190	12688
x"00",	-- Hex Addr	3191	12689
x"00",	-- Hex Addr	3192	12690
x"00",	-- Hex Addr	3193	12691
x"00",	-- Hex Addr	3194	12692
x"00",	-- Hex Addr	3195	12693
x"00",	-- Hex Addr	3196	12694
x"00",	-- Hex Addr	3197	12695
x"00",	-- Hex Addr	3198	12696
x"00",	-- Hex Addr	3199	12697
x"00",	-- Hex Addr	319A	12698
x"00",	-- Hex Addr	319B	12699
x"00",	-- Hex Addr	319C	12700
x"00",	-- Hex Addr	319D	12701
x"00",	-- Hex Addr	319E	12702
x"00",	-- Hex Addr	319F	12703
x"00",	-- Hex Addr	31A0	12704
x"00",	-- Hex Addr	31A1	12705
x"00",	-- Hex Addr	31A2	12706
x"00",	-- Hex Addr	31A3	12707
x"00",	-- Hex Addr	31A4	12708
x"00",	-- Hex Addr	31A5	12709
x"00",	-- Hex Addr	31A6	12710
x"00",	-- Hex Addr	31A7	12711
x"00",	-- Hex Addr	31A8	12712
x"00",	-- Hex Addr	31A9	12713
x"00",	-- Hex Addr	31AA	12714
x"00",	-- Hex Addr	31AB	12715
x"00",	-- Hex Addr	31AC	12716
x"00",	-- Hex Addr	31AD	12717
x"00",	-- Hex Addr	31AE	12718
x"00",	-- Hex Addr	31AF	12719
x"00",	-- Hex Addr	31B0	12720
x"00",	-- Hex Addr	31B1	12721
x"00",	-- Hex Addr	31B2	12722
x"00",	-- Hex Addr	31B3	12723
x"00",	-- Hex Addr	31B4	12724
x"00",	-- Hex Addr	31B5	12725
x"00",	-- Hex Addr	31B6	12726
x"00",	-- Hex Addr	31B7	12727
x"00",	-- Hex Addr	31B8	12728
x"00",	-- Hex Addr	31B9	12729
x"00",	-- Hex Addr	31BA	12730
x"00",	-- Hex Addr	31BB	12731
x"00",	-- Hex Addr	31BC	12732
x"00",	-- Hex Addr	31BD	12733
x"00",	-- Hex Addr	31BE	12734
x"00",	-- Hex Addr	31BF	12735
x"00",	-- Hex Addr	31C0	12736
x"00",	-- Hex Addr	31C1	12737
x"00",	-- Hex Addr	31C2	12738
x"00",	-- Hex Addr	31C3	12739
x"00",	-- Hex Addr	31C4	12740
x"00",	-- Hex Addr	31C5	12741
x"00",	-- Hex Addr	31C6	12742
x"00",	-- Hex Addr	31C7	12743
x"00",	-- Hex Addr	31C8	12744
x"00",	-- Hex Addr	31C9	12745
x"00",	-- Hex Addr	31CA	12746
x"00",	-- Hex Addr	31CB	12747
x"00",	-- Hex Addr	31CC	12748
x"00",	-- Hex Addr	31CD	12749
x"00",	-- Hex Addr	31CE	12750
x"00",	-- Hex Addr	31CF	12751
x"00",	-- Hex Addr	31D0	12752
x"00",	-- Hex Addr	31D1	12753
x"00",	-- Hex Addr	31D2	12754
x"00",	-- Hex Addr	31D3	12755
x"00",	-- Hex Addr	31D4	12756
x"00",	-- Hex Addr	31D5	12757
x"00",	-- Hex Addr	31D6	12758
x"00",	-- Hex Addr	31D7	12759
x"00",	-- Hex Addr	31D8	12760
x"00",	-- Hex Addr	31D9	12761
x"00",	-- Hex Addr	31DA	12762
x"00",	-- Hex Addr	31DB	12763
x"00",	-- Hex Addr	31DC	12764
x"00",	-- Hex Addr	31DD	12765
x"00",	-- Hex Addr	31DE	12766
x"00",	-- Hex Addr	31DF	12767
x"00",	-- Hex Addr	31E0	12768
x"00",	-- Hex Addr	31E1	12769
x"00",	-- Hex Addr	31E2	12770
x"00",	-- Hex Addr	31E3	12771
x"00",	-- Hex Addr	31E4	12772
x"00",	-- Hex Addr	31E5	12773
x"00",	-- Hex Addr	31E6	12774
x"00",	-- Hex Addr	31E7	12775
x"00",	-- Hex Addr	31E8	12776
x"00",	-- Hex Addr	31E9	12777
x"00",	-- Hex Addr	31EA	12778
x"00",	-- Hex Addr	31EB	12779
x"00",	-- Hex Addr	31EC	12780
x"00",	-- Hex Addr	31ED	12781
x"00",	-- Hex Addr	31EE	12782
x"00",	-- Hex Addr	31EF	12783
x"00",	-- Hex Addr	31F0	12784
x"00",	-- Hex Addr	31F1	12785
x"00",	-- Hex Addr	31F2	12786
x"00",	-- Hex Addr	31F3	12787
x"00",	-- Hex Addr	31F4	12788
x"00",	-- Hex Addr	31F5	12789
x"00",	-- Hex Addr	31F6	12790
x"00",	-- Hex Addr	31F7	12791
x"00",	-- Hex Addr	31F8	12792
x"00",	-- Hex Addr	31F9	12793
x"00",	-- Hex Addr	31FA	12794
x"00",	-- Hex Addr	31FB	12795
x"00",	-- Hex Addr	31FC	12796
x"00",	-- Hex Addr	31FD	12797
x"00",	-- Hex Addr	31FE	12798
x"00",	-- Hex Addr	31FF	12799
x"00",	-- Hex Addr	3200	12800
x"00",	-- Hex Addr	3201	12801
x"00",	-- Hex Addr	3202	12802
x"00",	-- Hex Addr	3203	12803
x"00",	-- Hex Addr	3204	12804
x"00",	-- Hex Addr	3205	12805
x"00",	-- Hex Addr	3206	12806
x"00",	-- Hex Addr	3207	12807
x"00",	-- Hex Addr	3208	12808
x"00",	-- Hex Addr	3209	12809
x"00",	-- Hex Addr	320A	12810
x"00",	-- Hex Addr	320B	12811
x"00",	-- Hex Addr	320C	12812
x"00",	-- Hex Addr	320D	12813
x"00",	-- Hex Addr	320E	12814
x"00",	-- Hex Addr	320F	12815
x"00",	-- Hex Addr	3210	12816
x"00",	-- Hex Addr	3211	12817
x"00",	-- Hex Addr	3212	12818
x"00",	-- Hex Addr	3213	12819
x"00",	-- Hex Addr	3214	12820
x"00",	-- Hex Addr	3215	12821
x"00",	-- Hex Addr	3216	12822
x"00",	-- Hex Addr	3217	12823
x"00",	-- Hex Addr	3218	12824
x"00",	-- Hex Addr	3219	12825
x"00",	-- Hex Addr	321A	12826
x"00",	-- Hex Addr	321B	12827
x"00",	-- Hex Addr	321C	12828
x"00",	-- Hex Addr	321D	12829
x"00",	-- Hex Addr	321E	12830
x"00",	-- Hex Addr	321F	12831
x"00",	-- Hex Addr	3220	12832
x"00",	-- Hex Addr	3221	12833
x"00",	-- Hex Addr	3222	12834
x"00",	-- Hex Addr	3223	12835
x"00",	-- Hex Addr	3224	12836
x"00",	-- Hex Addr	3225	12837
x"00",	-- Hex Addr	3226	12838
x"00",	-- Hex Addr	3227	12839
x"00",	-- Hex Addr	3228	12840
x"00",	-- Hex Addr	3229	12841
x"00",	-- Hex Addr	322A	12842
x"00",	-- Hex Addr	322B	12843
x"00",	-- Hex Addr	322C	12844
x"00",	-- Hex Addr	322D	12845
x"00",	-- Hex Addr	322E	12846
x"00",	-- Hex Addr	322F	12847
x"00",	-- Hex Addr	3230	12848
x"00",	-- Hex Addr	3231	12849
x"00",	-- Hex Addr	3232	12850
x"00",	-- Hex Addr	3233	12851
x"00",	-- Hex Addr	3234	12852
x"00",	-- Hex Addr	3235	12853
x"00",	-- Hex Addr	3236	12854
x"00",	-- Hex Addr	3237	12855
x"00",	-- Hex Addr	3238	12856
x"00",	-- Hex Addr	3239	12857
x"00",	-- Hex Addr	323A	12858
x"00",	-- Hex Addr	323B	12859
x"00",	-- Hex Addr	323C	12860
x"00",	-- Hex Addr	323D	12861
x"00",	-- Hex Addr	323E	12862
x"00",	-- Hex Addr	323F	12863
x"00",	-- Hex Addr	3240	12864
x"00",	-- Hex Addr	3241	12865
x"00",	-- Hex Addr	3242	12866
x"00",	-- Hex Addr	3243	12867
x"00",	-- Hex Addr	3244	12868
x"00",	-- Hex Addr	3245	12869
x"00",	-- Hex Addr	3246	12870
x"00",	-- Hex Addr	3247	12871
x"00",	-- Hex Addr	3248	12872
x"00",	-- Hex Addr	3249	12873
x"00",	-- Hex Addr	324A	12874
x"00",	-- Hex Addr	324B	12875
x"00",	-- Hex Addr	324C	12876
x"00",	-- Hex Addr	324D	12877
x"00",	-- Hex Addr	324E	12878
x"00",	-- Hex Addr	324F	12879
x"00",	-- Hex Addr	3250	12880
x"00",	-- Hex Addr	3251	12881
x"00",	-- Hex Addr	3252	12882
x"00",	-- Hex Addr	3253	12883
x"00",	-- Hex Addr	3254	12884
x"00",	-- Hex Addr	3255	12885
x"00",	-- Hex Addr	3256	12886
x"00",	-- Hex Addr	3257	12887
x"00",	-- Hex Addr	3258	12888
x"00",	-- Hex Addr	3259	12889
x"00",	-- Hex Addr	325A	12890
x"00",	-- Hex Addr	325B	12891
x"00",	-- Hex Addr	325C	12892
x"00",	-- Hex Addr	325D	12893
x"00",	-- Hex Addr	325E	12894
x"00",	-- Hex Addr	325F	12895
x"00",	-- Hex Addr	3260	12896
x"00",	-- Hex Addr	3261	12897
x"00",	-- Hex Addr	3262	12898
x"00",	-- Hex Addr	3263	12899
x"00",	-- Hex Addr	3264	12900
x"00",	-- Hex Addr	3265	12901
x"00",	-- Hex Addr	3266	12902
x"00",	-- Hex Addr	3267	12903
x"00",	-- Hex Addr	3268	12904
x"00",	-- Hex Addr	3269	12905
x"00",	-- Hex Addr	326A	12906
x"00",	-- Hex Addr	326B	12907
x"00",	-- Hex Addr	326C	12908
x"00",	-- Hex Addr	326D	12909
x"00",	-- Hex Addr	326E	12910
x"00",	-- Hex Addr	326F	12911
x"00",	-- Hex Addr	3270	12912
x"00",	-- Hex Addr	3271	12913
x"00",	-- Hex Addr	3272	12914
x"00",	-- Hex Addr	3273	12915
x"00",	-- Hex Addr	3274	12916
x"00",	-- Hex Addr	3275	12917
x"00",	-- Hex Addr	3276	12918
x"00",	-- Hex Addr	3277	12919
x"00",	-- Hex Addr	3278	12920
x"00",	-- Hex Addr	3279	12921
x"00",	-- Hex Addr	327A	12922
x"00",	-- Hex Addr	327B	12923
x"00",	-- Hex Addr	327C	12924
x"00",	-- Hex Addr	327D	12925
x"00",	-- Hex Addr	327E	12926
x"00",	-- Hex Addr	327F	12927
x"00",	-- Hex Addr	3280	12928
x"00",	-- Hex Addr	3281	12929
x"00",	-- Hex Addr	3282	12930
x"00",	-- Hex Addr	3283	12931
x"00",	-- Hex Addr	3284	12932
x"00",	-- Hex Addr	3285	12933
x"00",	-- Hex Addr	3286	12934
x"00",	-- Hex Addr	3287	12935
x"00",	-- Hex Addr	3288	12936
x"00",	-- Hex Addr	3289	12937
x"00",	-- Hex Addr	328A	12938
x"00",	-- Hex Addr	328B	12939
x"00",	-- Hex Addr	328C	12940
x"00",	-- Hex Addr	328D	12941
x"00",	-- Hex Addr	328E	12942
x"00",	-- Hex Addr	328F	12943
x"00",	-- Hex Addr	3290	12944
x"00",	-- Hex Addr	3291	12945
x"00",	-- Hex Addr	3292	12946
x"00",	-- Hex Addr	3293	12947
x"00",	-- Hex Addr	3294	12948
x"00",	-- Hex Addr	3295	12949
x"00",	-- Hex Addr	3296	12950
x"00",	-- Hex Addr	3297	12951
x"00",	-- Hex Addr	3298	12952
x"00",	-- Hex Addr	3299	12953
x"00",	-- Hex Addr	329A	12954
x"00",	-- Hex Addr	329B	12955
x"00",	-- Hex Addr	329C	12956
x"00",	-- Hex Addr	329D	12957
x"00",	-- Hex Addr	329E	12958
x"00",	-- Hex Addr	329F	12959
x"00",	-- Hex Addr	32A0	12960
x"00",	-- Hex Addr	32A1	12961
x"00",	-- Hex Addr	32A2	12962
x"00",	-- Hex Addr	32A3	12963
x"00",	-- Hex Addr	32A4	12964
x"00",	-- Hex Addr	32A5	12965
x"00",	-- Hex Addr	32A6	12966
x"00",	-- Hex Addr	32A7	12967
x"00",	-- Hex Addr	32A8	12968
x"00",	-- Hex Addr	32A9	12969
x"00",	-- Hex Addr	32AA	12970
x"00",	-- Hex Addr	32AB	12971
x"00",	-- Hex Addr	32AC	12972
x"00",	-- Hex Addr	32AD	12973
x"00",	-- Hex Addr	32AE	12974
x"00",	-- Hex Addr	32AF	12975
x"00",	-- Hex Addr	32B0	12976
x"00",	-- Hex Addr	32B1	12977
x"00",	-- Hex Addr	32B2	12978
x"00",	-- Hex Addr	32B3	12979
x"00",	-- Hex Addr	32B4	12980
x"00",	-- Hex Addr	32B5	12981
x"00",	-- Hex Addr	32B6	12982
x"00",	-- Hex Addr	32B7	12983
x"00",	-- Hex Addr	32B8	12984
x"00",	-- Hex Addr	32B9	12985
x"00",	-- Hex Addr	32BA	12986
x"00",	-- Hex Addr	32BB	12987
x"00",	-- Hex Addr	32BC	12988
x"00",	-- Hex Addr	32BD	12989
x"00",	-- Hex Addr	32BE	12990
x"00",	-- Hex Addr	32BF	12991
x"00",	-- Hex Addr	32C0	12992
x"00",	-- Hex Addr	32C1	12993
x"00",	-- Hex Addr	32C2	12994
x"00",	-- Hex Addr	32C3	12995
x"00",	-- Hex Addr	32C4	12996
x"00",	-- Hex Addr	32C5	12997
x"00",	-- Hex Addr	32C6	12998
x"00",	-- Hex Addr	32C7	12999
x"00",	-- Hex Addr	32C8	13000
x"00",	-- Hex Addr	32C9	13001
x"00",	-- Hex Addr	32CA	13002
x"00",	-- Hex Addr	32CB	13003
x"00",	-- Hex Addr	32CC	13004
x"00",	-- Hex Addr	32CD	13005
x"00",	-- Hex Addr	32CE	13006
x"00",	-- Hex Addr	32CF	13007
x"00",	-- Hex Addr	32D0	13008
x"00",	-- Hex Addr	32D1	13009
x"00",	-- Hex Addr	32D2	13010
x"00",	-- Hex Addr	32D3	13011
x"00",	-- Hex Addr	32D4	13012
x"00",	-- Hex Addr	32D5	13013
x"00",	-- Hex Addr	32D6	13014
x"00",	-- Hex Addr	32D7	13015
x"00",	-- Hex Addr	32D8	13016
x"00",	-- Hex Addr	32D9	13017
x"00",	-- Hex Addr	32DA	13018
x"00",	-- Hex Addr	32DB	13019
x"00",	-- Hex Addr	32DC	13020
x"00",	-- Hex Addr	32DD	13021
x"00",	-- Hex Addr	32DE	13022
x"00",	-- Hex Addr	32DF	13023
x"00",	-- Hex Addr	32E0	13024
x"00",	-- Hex Addr	32E1	13025
x"00",	-- Hex Addr	32E2	13026
x"00",	-- Hex Addr	32E3	13027
x"00",	-- Hex Addr	32E4	13028
x"00",	-- Hex Addr	32E5	13029
x"00",	-- Hex Addr	32E6	13030
x"00",	-- Hex Addr	32E7	13031
x"00",	-- Hex Addr	32E8	13032
x"00",	-- Hex Addr	32E9	13033
x"00",	-- Hex Addr	32EA	13034
x"00",	-- Hex Addr	32EB	13035
x"00",	-- Hex Addr	32EC	13036
x"00",	-- Hex Addr	32ED	13037
x"00",	-- Hex Addr	32EE	13038
x"00",	-- Hex Addr	32EF	13039
x"00",	-- Hex Addr	32F0	13040
x"00",	-- Hex Addr	32F1	13041
x"00",	-- Hex Addr	32F2	13042
x"00",	-- Hex Addr	32F3	13043
x"00",	-- Hex Addr	32F4	13044
x"00",	-- Hex Addr	32F5	13045
x"00",	-- Hex Addr	32F6	13046
x"00",	-- Hex Addr	32F7	13047
x"00",	-- Hex Addr	32F8	13048
x"00",	-- Hex Addr	32F9	13049
x"00",	-- Hex Addr	32FA	13050
x"00",	-- Hex Addr	32FB	13051
x"00",	-- Hex Addr	32FC	13052
x"00",	-- Hex Addr	32FD	13053
x"00",	-- Hex Addr	32FE	13054
x"00",	-- Hex Addr	32FF	13055
x"00",	-- Hex Addr	3300	13056
x"00",	-- Hex Addr	3301	13057
x"00",	-- Hex Addr	3302	13058
x"00",	-- Hex Addr	3303	13059
x"00",	-- Hex Addr	3304	13060
x"00",	-- Hex Addr	3305	13061
x"00",	-- Hex Addr	3306	13062
x"00",	-- Hex Addr	3307	13063
x"00",	-- Hex Addr	3308	13064
x"00",	-- Hex Addr	3309	13065
x"00",	-- Hex Addr	330A	13066
x"00",	-- Hex Addr	330B	13067
x"00",	-- Hex Addr	330C	13068
x"00",	-- Hex Addr	330D	13069
x"00",	-- Hex Addr	330E	13070
x"00",	-- Hex Addr	330F	13071
x"00",	-- Hex Addr	3310	13072
x"00",	-- Hex Addr	3311	13073
x"00",	-- Hex Addr	3312	13074
x"00",	-- Hex Addr	3313	13075
x"00",	-- Hex Addr	3314	13076
x"00",	-- Hex Addr	3315	13077
x"00",	-- Hex Addr	3316	13078
x"00",	-- Hex Addr	3317	13079
x"00",	-- Hex Addr	3318	13080
x"00",	-- Hex Addr	3319	13081
x"00",	-- Hex Addr	331A	13082
x"00",	-- Hex Addr	331B	13083
x"00",	-- Hex Addr	331C	13084
x"00",	-- Hex Addr	331D	13085
x"00",	-- Hex Addr	331E	13086
x"00",	-- Hex Addr	331F	13087
x"00",	-- Hex Addr	3320	13088
x"00",	-- Hex Addr	3321	13089
x"00",	-- Hex Addr	3322	13090
x"00",	-- Hex Addr	3323	13091
x"00",	-- Hex Addr	3324	13092
x"00",	-- Hex Addr	3325	13093
x"00",	-- Hex Addr	3326	13094
x"00",	-- Hex Addr	3327	13095
x"00",	-- Hex Addr	3328	13096
x"00",	-- Hex Addr	3329	13097
x"00",	-- Hex Addr	332A	13098
x"00",	-- Hex Addr	332B	13099
x"00",	-- Hex Addr	332C	13100
x"00",	-- Hex Addr	332D	13101
x"00",	-- Hex Addr	332E	13102
x"00",	-- Hex Addr	332F	13103
x"00",	-- Hex Addr	3330	13104
x"00",	-- Hex Addr	3331	13105
x"00",	-- Hex Addr	3332	13106
x"00",	-- Hex Addr	3333	13107
x"00",	-- Hex Addr	3334	13108
x"00",	-- Hex Addr	3335	13109
x"00",	-- Hex Addr	3336	13110
x"00",	-- Hex Addr	3337	13111
x"00",	-- Hex Addr	3338	13112
x"00",	-- Hex Addr	3339	13113
x"00",	-- Hex Addr	333A	13114
x"00",	-- Hex Addr	333B	13115
x"00",	-- Hex Addr	333C	13116
x"00",	-- Hex Addr	333D	13117
x"00",	-- Hex Addr	333E	13118
x"00",	-- Hex Addr	333F	13119
x"00",	-- Hex Addr	3340	13120
x"00",	-- Hex Addr	3341	13121
x"00",	-- Hex Addr	3342	13122
x"00",	-- Hex Addr	3343	13123
x"00",	-- Hex Addr	3344	13124
x"00",	-- Hex Addr	3345	13125
x"00",	-- Hex Addr	3346	13126
x"00",	-- Hex Addr	3347	13127
x"00",	-- Hex Addr	3348	13128
x"00",	-- Hex Addr	3349	13129
x"00",	-- Hex Addr	334A	13130
x"00",	-- Hex Addr	334B	13131
x"00",	-- Hex Addr	334C	13132
x"00",	-- Hex Addr	334D	13133
x"00",	-- Hex Addr	334E	13134
x"00",	-- Hex Addr	334F	13135
x"00",	-- Hex Addr	3350	13136
x"00",	-- Hex Addr	3351	13137
x"00",	-- Hex Addr	3352	13138
x"00",	-- Hex Addr	3353	13139
x"00",	-- Hex Addr	3354	13140
x"00",	-- Hex Addr	3355	13141
x"00",	-- Hex Addr	3356	13142
x"00",	-- Hex Addr	3357	13143
x"00",	-- Hex Addr	3358	13144
x"00",	-- Hex Addr	3359	13145
x"00",	-- Hex Addr	335A	13146
x"00",	-- Hex Addr	335B	13147
x"00",	-- Hex Addr	335C	13148
x"00",	-- Hex Addr	335D	13149
x"00",	-- Hex Addr	335E	13150
x"00",	-- Hex Addr	335F	13151
x"00",	-- Hex Addr	3360	13152
x"00",	-- Hex Addr	3361	13153
x"00",	-- Hex Addr	3362	13154
x"00",	-- Hex Addr	3363	13155
x"00",	-- Hex Addr	3364	13156
x"00",	-- Hex Addr	3365	13157
x"00",	-- Hex Addr	3366	13158
x"00",	-- Hex Addr	3367	13159
x"00",	-- Hex Addr	3368	13160
x"00",	-- Hex Addr	3369	13161
x"00",	-- Hex Addr	336A	13162
x"00",	-- Hex Addr	336B	13163
x"00",	-- Hex Addr	336C	13164
x"00",	-- Hex Addr	336D	13165
x"00",	-- Hex Addr	336E	13166
x"00",	-- Hex Addr	336F	13167
x"00",	-- Hex Addr	3370	13168
x"00",	-- Hex Addr	3371	13169
x"00",	-- Hex Addr	3372	13170
x"00",	-- Hex Addr	3373	13171
x"00",	-- Hex Addr	3374	13172
x"00",	-- Hex Addr	3375	13173
x"00",	-- Hex Addr	3376	13174
x"00",	-- Hex Addr	3377	13175
x"00",	-- Hex Addr	3378	13176
x"00",	-- Hex Addr	3379	13177
x"00",	-- Hex Addr	337A	13178
x"00",	-- Hex Addr	337B	13179
x"00",	-- Hex Addr	337C	13180
x"00",	-- Hex Addr	337D	13181
x"00",	-- Hex Addr	337E	13182
x"00",	-- Hex Addr	337F	13183
x"00",	-- Hex Addr	3380	13184
x"00",	-- Hex Addr	3381	13185
x"00",	-- Hex Addr	3382	13186
x"00",	-- Hex Addr	3383	13187
x"00",	-- Hex Addr	3384	13188
x"00",	-- Hex Addr	3385	13189
x"00",	-- Hex Addr	3386	13190
x"00",	-- Hex Addr	3387	13191
x"00",	-- Hex Addr	3388	13192
x"00",	-- Hex Addr	3389	13193
x"00",	-- Hex Addr	338A	13194
x"00",	-- Hex Addr	338B	13195
x"00",	-- Hex Addr	338C	13196
x"00",	-- Hex Addr	338D	13197
x"00",	-- Hex Addr	338E	13198
x"00",	-- Hex Addr	338F	13199
x"00",	-- Hex Addr	3390	13200
x"00",	-- Hex Addr	3391	13201
x"00",	-- Hex Addr	3392	13202
x"00",	-- Hex Addr	3393	13203
x"00",	-- Hex Addr	3394	13204
x"00",	-- Hex Addr	3395	13205
x"00",	-- Hex Addr	3396	13206
x"00",	-- Hex Addr	3397	13207
x"00",	-- Hex Addr	3398	13208
x"00",	-- Hex Addr	3399	13209
x"00",	-- Hex Addr	339A	13210
x"00",	-- Hex Addr	339B	13211
x"00",	-- Hex Addr	339C	13212
x"00",	-- Hex Addr	339D	13213
x"00",	-- Hex Addr	339E	13214
x"00",	-- Hex Addr	339F	13215
x"00",	-- Hex Addr	33A0	13216
x"00",	-- Hex Addr	33A1	13217
x"00",	-- Hex Addr	33A2	13218
x"00",	-- Hex Addr	33A3	13219
x"00",	-- Hex Addr	33A4	13220
x"00",	-- Hex Addr	33A5	13221
x"00",	-- Hex Addr	33A6	13222
x"00",	-- Hex Addr	33A7	13223
x"00",	-- Hex Addr	33A8	13224
x"00",	-- Hex Addr	33A9	13225
x"00",	-- Hex Addr	33AA	13226
x"00",	-- Hex Addr	33AB	13227
x"00",	-- Hex Addr	33AC	13228
x"00",	-- Hex Addr	33AD	13229
x"00",	-- Hex Addr	33AE	13230
x"00",	-- Hex Addr	33AF	13231
x"00",	-- Hex Addr	33B0	13232
x"00",	-- Hex Addr	33B1	13233
x"00",	-- Hex Addr	33B2	13234
x"00",	-- Hex Addr	33B3	13235
x"00",	-- Hex Addr	33B4	13236
x"00",	-- Hex Addr	33B5	13237
x"00",	-- Hex Addr	33B6	13238
x"00",	-- Hex Addr	33B7	13239
x"00",	-- Hex Addr	33B8	13240
x"00",	-- Hex Addr	33B9	13241
x"00",	-- Hex Addr	33BA	13242
x"00",	-- Hex Addr	33BB	13243
x"00",	-- Hex Addr	33BC	13244
x"00",	-- Hex Addr	33BD	13245
x"00",	-- Hex Addr	33BE	13246
x"00",	-- Hex Addr	33BF	13247
x"00",	-- Hex Addr	33C0	13248
x"00",	-- Hex Addr	33C1	13249
x"00",	-- Hex Addr	33C2	13250
x"00",	-- Hex Addr	33C3	13251
x"00",	-- Hex Addr	33C4	13252
x"00",	-- Hex Addr	33C5	13253
x"00",	-- Hex Addr	33C6	13254
x"00",	-- Hex Addr	33C7	13255
x"00",	-- Hex Addr	33C8	13256
x"00",	-- Hex Addr	33C9	13257
x"00",	-- Hex Addr	33CA	13258
x"00",	-- Hex Addr	33CB	13259
x"00",	-- Hex Addr	33CC	13260
x"00",	-- Hex Addr	33CD	13261
x"00",	-- Hex Addr	33CE	13262
x"00",	-- Hex Addr	33CF	13263
x"00",	-- Hex Addr	33D0	13264
x"00",	-- Hex Addr	33D1	13265
x"00",	-- Hex Addr	33D2	13266
x"00",	-- Hex Addr	33D3	13267
x"00",	-- Hex Addr	33D4	13268
x"00",	-- Hex Addr	33D5	13269
x"00",	-- Hex Addr	33D6	13270
x"00",	-- Hex Addr	33D7	13271
x"00",	-- Hex Addr	33D8	13272
x"00",	-- Hex Addr	33D9	13273
x"00",	-- Hex Addr	33DA	13274
x"00",	-- Hex Addr	33DB	13275
x"00",	-- Hex Addr	33DC	13276
x"00",	-- Hex Addr	33DD	13277
x"00",	-- Hex Addr	33DE	13278
x"00",	-- Hex Addr	33DF	13279
x"00",	-- Hex Addr	33E0	13280
x"00",	-- Hex Addr	33E1	13281
x"00",	-- Hex Addr	33E2	13282
x"00",	-- Hex Addr	33E3	13283
x"00",	-- Hex Addr	33E4	13284
x"00",	-- Hex Addr	33E5	13285
x"00",	-- Hex Addr	33E6	13286
x"00",	-- Hex Addr	33E7	13287
x"00",	-- Hex Addr	33E8	13288
x"00",	-- Hex Addr	33E9	13289
x"00",	-- Hex Addr	33EA	13290
x"00",	-- Hex Addr	33EB	13291
x"00",	-- Hex Addr	33EC	13292
x"00",	-- Hex Addr	33ED	13293
x"00",	-- Hex Addr	33EE	13294
x"00",	-- Hex Addr	33EF	13295
x"00",	-- Hex Addr	33F0	13296
x"00",	-- Hex Addr	33F1	13297
x"00",	-- Hex Addr	33F2	13298
x"00",	-- Hex Addr	33F3	13299
x"00",	-- Hex Addr	33F4	13300
x"00",	-- Hex Addr	33F5	13301
x"00",	-- Hex Addr	33F6	13302
x"00",	-- Hex Addr	33F7	13303
x"00",	-- Hex Addr	33F8	13304
x"00",	-- Hex Addr	33F9	13305
x"00",	-- Hex Addr	33FA	13306
x"00",	-- Hex Addr	33FB	13307
x"00",	-- Hex Addr	33FC	13308
x"00",	-- Hex Addr	33FD	13309
x"00",	-- Hex Addr	33FE	13310
x"00",	-- Hex Addr	33FF	13311
x"00",	-- Hex Addr	3400	13312
x"00",	-- Hex Addr	3401	13313
x"00",	-- Hex Addr	3402	13314
x"00",	-- Hex Addr	3403	13315
x"00",	-- Hex Addr	3404	13316
x"00",	-- Hex Addr	3405	13317
x"00",	-- Hex Addr	3406	13318
x"00",	-- Hex Addr	3407	13319
x"00",	-- Hex Addr	3408	13320
x"00",	-- Hex Addr	3409	13321
x"00",	-- Hex Addr	340A	13322
x"00",	-- Hex Addr	340B	13323
x"00",	-- Hex Addr	340C	13324
x"00",	-- Hex Addr	340D	13325
x"00",	-- Hex Addr	340E	13326
x"00",	-- Hex Addr	340F	13327
x"00",	-- Hex Addr	3410	13328
x"00",	-- Hex Addr	3411	13329
x"00",	-- Hex Addr	3412	13330
x"00",	-- Hex Addr	3413	13331
x"00",	-- Hex Addr	3414	13332
x"00",	-- Hex Addr	3415	13333
x"00",	-- Hex Addr	3416	13334
x"00",	-- Hex Addr	3417	13335
x"00",	-- Hex Addr	3418	13336
x"00",	-- Hex Addr	3419	13337
x"00",	-- Hex Addr	341A	13338
x"00",	-- Hex Addr	341B	13339
x"00",	-- Hex Addr	341C	13340
x"00",	-- Hex Addr	341D	13341
x"00",	-- Hex Addr	341E	13342
x"00",	-- Hex Addr	341F	13343
x"00",	-- Hex Addr	3420	13344
x"00",	-- Hex Addr	3421	13345
x"00",	-- Hex Addr	3422	13346
x"00",	-- Hex Addr	3423	13347
x"00",	-- Hex Addr	3424	13348
x"00",	-- Hex Addr	3425	13349
x"00",	-- Hex Addr	3426	13350
x"00",	-- Hex Addr	3427	13351
x"00",	-- Hex Addr	3428	13352
x"00",	-- Hex Addr	3429	13353
x"00",	-- Hex Addr	342A	13354
x"00",	-- Hex Addr	342B	13355
x"00",	-- Hex Addr	342C	13356
x"00",	-- Hex Addr	342D	13357
x"00",	-- Hex Addr	342E	13358
x"00",	-- Hex Addr	342F	13359
x"00",	-- Hex Addr	3430	13360
x"00",	-- Hex Addr	3431	13361
x"00",	-- Hex Addr	3432	13362
x"00",	-- Hex Addr	3433	13363
x"00",	-- Hex Addr	3434	13364
x"00",	-- Hex Addr	3435	13365
x"00",	-- Hex Addr	3436	13366
x"00",	-- Hex Addr	3437	13367
x"00",	-- Hex Addr	3438	13368
x"00",	-- Hex Addr	3439	13369
x"00",	-- Hex Addr	343A	13370
x"00",	-- Hex Addr	343B	13371
x"00",	-- Hex Addr	343C	13372
x"00",	-- Hex Addr	343D	13373
x"00",	-- Hex Addr	343E	13374
x"00",	-- Hex Addr	343F	13375
x"00",	-- Hex Addr	3440	13376
x"00",	-- Hex Addr	3441	13377
x"00",	-- Hex Addr	3442	13378
x"00",	-- Hex Addr	3443	13379
x"00",	-- Hex Addr	3444	13380
x"00",	-- Hex Addr	3445	13381
x"00",	-- Hex Addr	3446	13382
x"00",	-- Hex Addr	3447	13383
x"00",	-- Hex Addr	3448	13384
x"00",	-- Hex Addr	3449	13385
x"00",	-- Hex Addr	344A	13386
x"00",	-- Hex Addr	344B	13387
x"00",	-- Hex Addr	344C	13388
x"00",	-- Hex Addr	344D	13389
x"00",	-- Hex Addr	344E	13390
x"00",	-- Hex Addr	344F	13391
x"00",	-- Hex Addr	3450	13392
x"00",	-- Hex Addr	3451	13393
x"00",	-- Hex Addr	3452	13394
x"00",	-- Hex Addr	3453	13395
x"00",	-- Hex Addr	3454	13396
x"00",	-- Hex Addr	3455	13397
x"00",	-- Hex Addr	3456	13398
x"00",	-- Hex Addr	3457	13399
x"00",	-- Hex Addr	3458	13400
x"00",	-- Hex Addr	3459	13401
x"00",	-- Hex Addr	345A	13402
x"00",	-- Hex Addr	345B	13403
x"00",	-- Hex Addr	345C	13404
x"00",	-- Hex Addr	345D	13405
x"00",	-- Hex Addr	345E	13406
x"00",	-- Hex Addr	345F	13407
x"00",	-- Hex Addr	3460	13408
x"00",	-- Hex Addr	3461	13409
x"00",	-- Hex Addr	3462	13410
x"00",	-- Hex Addr	3463	13411
x"00",	-- Hex Addr	3464	13412
x"00",	-- Hex Addr	3465	13413
x"00",	-- Hex Addr	3466	13414
x"00",	-- Hex Addr	3467	13415
x"00",	-- Hex Addr	3468	13416
x"00",	-- Hex Addr	3469	13417
x"00",	-- Hex Addr	346A	13418
x"00",	-- Hex Addr	346B	13419
x"00",	-- Hex Addr	346C	13420
x"00",	-- Hex Addr	346D	13421
x"00",	-- Hex Addr	346E	13422
x"00",	-- Hex Addr	346F	13423
x"00",	-- Hex Addr	3470	13424
x"00",	-- Hex Addr	3471	13425
x"00",	-- Hex Addr	3472	13426
x"00",	-- Hex Addr	3473	13427
x"00",	-- Hex Addr	3474	13428
x"00",	-- Hex Addr	3475	13429
x"00",	-- Hex Addr	3476	13430
x"00",	-- Hex Addr	3477	13431
x"00",	-- Hex Addr	3478	13432
x"00",	-- Hex Addr	3479	13433
x"00",	-- Hex Addr	347A	13434
x"00",	-- Hex Addr	347B	13435
x"00",	-- Hex Addr	347C	13436
x"00",	-- Hex Addr	347D	13437
x"00",	-- Hex Addr	347E	13438
x"00",	-- Hex Addr	347F	13439
x"00",	-- Hex Addr	3480	13440
x"00",	-- Hex Addr	3481	13441
x"00",	-- Hex Addr	3482	13442
x"00",	-- Hex Addr	3483	13443
x"00",	-- Hex Addr	3484	13444
x"00",	-- Hex Addr	3485	13445
x"00",	-- Hex Addr	3486	13446
x"00",	-- Hex Addr	3487	13447
x"00",	-- Hex Addr	3488	13448
x"00",	-- Hex Addr	3489	13449
x"00",	-- Hex Addr	348A	13450
x"00",	-- Hex Addr	348B	13451
x"00",	-- Hex Addr	348C	13452
x"00",	-- Hex Addr	348D	13453
x"00",	-- Hex Addr	348E	13454
x"00",	-- Hex Addr	348F	13455
x"00",	-- Hex Addr	3490	13456
x"00",	-- Hex Addr	3491	13457
x"00",	-- Hex Addr	3492	13458
x"00",	-- Hex Addr	3493	13459
x"00",	-- Hex Addr	3494	13460
x"00",	-- Hex Addr	3495	13461
x"00",	-- Hex Addr	3496	13462
x"00",	-- Hex Addr	3497	13463
x"00",	-- Hex Addr	3498	13464
x"00",	-- Hex Addr	3499	13465
x"00",	-- Hex Addr	349A	13466
x"00",	-- Hex Addr	349B	13467
x"00",	-- Hex Addr	349C	13468
x"00",	-- Hex Addr	349D	13469
x"00",	-- Hex Addr	349E	13470
x"00",	-- Hex Addr	349F	13471
x"00",	-- Hex Addr	34A0	13472
x"00",	-- Hex Addr	34A1	13473
x"00",	-- Hex Addr	34A2	13474
x"00",	-- Hex Addr	34A3	13475
x"00",	-- Hex Addr	34A4	13476
x"00",	-- Hex Addr	34A5	13477
x"00",	-- Hex Addr	34A6	13478
x"00",	-- Hex Addr	34A7	13479
x"00",	-- Hex Addr	34A8	13480
x"00",	-- Hex Addr	34A9	13481
x"00",	-- Hex Addr	34AA	13482
x"00",	-- Hex Addr	34AB	13483
x"00",	-- Hex Addr	34AC	13484
x"00",	-- Hex Addr	34AD	13485
x"00",	-- Hex Addr	34AE	13486
x"00",	-- Hex Addr	34AF	13487
x"00",	-- Hex Addr	34B0	13488
x"00",	-- Hex Addr	34B1	13489
x"00",	-- Hex Addr	34B2	13490
x"00",	-- Hex Addr	34B3	13491
x"00",	-- Hex Addr	34B4	13492
x"00",	-- Hex Addr	34B5	13493
x"00",	-- Hex Addr	34B6	13494
x"00",	-- Hex Addr	34B7	13495
x"00",	-- Hex Addr	34B8	13496
x"00",	-- Hex Addr	34B9	13497
x"00",	-- Hex Addr	34BA	13498
x"00",	-- Hex Addr	34BB	13499
x"00",	-- Hex Addr	34BC	13500
x"00",	-- Hex Addr	34BD	13501
x"00",	-- Hex Addr	34BE	13502
x"00",	-- Hex Addr	34BF	13503
x"00",	-- Hex Addr	34C0	13504
x"00",	-- Hex Addr	34C1	13505
x"00",	-- Hex Addr	34C2	13506
x"00",	-- Hex Addr	34C3	13507
x"00",	-- Hex Addr	34C4	13508
x"00",	-- Hex Addr	34C5	13509
x"00",	-- Hex Addr	34C6	13510
x"00",	-- Hex Addr	34C7	13511
x"00",	-- Hex Addr	34C8	13512
x"00",	-- Hex Addr	34C9	13513
x"00",	-- Hex Addr	34CA	13514
x"00",	-- Hex Addr	34CB	13515
x"00",	-- Hex Addr	34CC	13516
x"00",	-- Hex Addr	34CD	13517
x"00",	-- Hex Addr	34CE	13518
x"00",	-- Hex Addr	34CF	13519
x"00",	-- Hex Addr	34D0	13520
x"00",	-- Hex Addr	34D1	13521
x"00",	-- Hex Addr	34D2	13522
x"00",	-- Hex Addr	34D3	13523
x"00",	-- Hex Addr	34D4	13524
x"00",	-- Hex Addr	34D5	13525
x"00",	-- Hex Addr	34D6	13526
x"00",	-- Hex Addr	34D7	13527
x"00",	-- Hex Addr	34D8	13528
x"00",	-- Hex Addr	34D9	13529
x"00",	-- Hex Addr	34DA	13530
x"00",	-- Hex Addr	34DB	13531
x"00",	-- Hex Addr	34DC	13532
x"00",	-- Hex Addr	34DD	13533
x"00",	-- Hex Addr	34DE	13534
x"00",	-- Hex Addr	34DF	13535
x"00",	-- Hex Addr	34E0	13536
x"00",	-- Hex Addr	34E1	13537
x"00",	-- Hex Addr	34E2	13538
x"00",	-- Hex Addr	34E3	13539
x"00",	-- Hex Addr	34E4	13540
x"00",	-- Hex Addr	34E5	13541
x"00",	-- Hex Addr	34E6	13542
x"00",	-- Hex Addr	34E7	13543
x"00",	-- Hex Addr	34E8	13544
x"00",	-- Hex Addr	34E9	13545
x"00",	-- Hex Addr	34EA	13546
x"00",	-- Hex Addr	34EB	13547
x"00",	-- Hex Addr	34EC	13548
x"00",	-- Hex Addr	34ED	13549
x"00",	-- Hex Addr	34EE	13550
x"00",	-- Hex Addr	34EF	13551
x"00",	-- Hex Addr	34F0	13552
x"00",	-- Hex Addr	34F1	13553
x"00",	-- Hex Addr	34F2	13554
x"00",	-- Hex Addr	34F3	13555
x"00",	-- Hex Addr	34F4	13556
x"00",	-- Hex Addr	34F5	13557
x"00",	-- Hex Addr	34F6	13558
x"00",	-- Hex Addr	34F7	13559
x"00",	-- Hex Addr	34F8	13560
x"00",	-- Hex Addr	34F9	13561
x"00",	-- Hex Addr	34FA	13562
x"00",	-- Hex Addr	34FB	13563
x"00",	-- Hex Addr	34FC	13564
x"00",	-- Hex Addr	34FD	13565
x"00",	-- Hex Addr	34FE	13566
x"00",	-- Hex Addr	34FF	13567
x"00",	-- Hex Addr	3500	13568
x"00",	-- Hex Addr	3501	13569
x"00",	-- Hex Addr	3502	13570
x"00",	-- Hex Addr	3503	13571
x"00",	-- Hex Addr	3504	13572
x"00",	-- Hex Addr	3505	13573
x"00",	-- Hex Addr	3506	13574
x"00",	-- Hex Addr	3507	13575
x"00",	-- Hex Addr	3508	13576
x"00",	-- Hex Addr	3509	13577
x"00",	-- Hex Addr	350A	13578
x"00",	-- Hex Addr	350B	13579
x"00",	-- Hex Addr	350C	13580
x"00",	-- Hex Addr	350D	13581
x"00",	-- Hex Addr	350E	13582
x"00",	-- Hex Addr	350F	13583
x"00",	-- Hex Addr	3510	13584
x"00",	-- Hex Addr	3511	13585
x"00",	-- Hex Addr	3512	13586
x"00",	-- Hex Addr	3513	13587
x"00",	-- Hex Addr	3514	13588
x"00",	-- Hex Addr	3515	13589
x"00",	-- Hex Addr	3516	13590
x"00",	-- Hex Addr	3517	13591
x"00",	-- Hex Addr	3518	13592
x"00",	-- Hex Addr	3519	13593
x"00",	-- Hex Addr	351A	13594
x"00",	-- Hex Addr	351B	13595
x"00",	-- Hex Addr	351C	13596
x"00",	-- Hex Addr	351D	13597
x"00",	-- Hex Addr	351E	13598
x"00",	-- Hex Addr	351F	13599
x"00",	-- Hex Addr	3520	13600
x"00",	-- Hex Addr	3521	13601
x"00",	-- Hex Addr	3522	13602
x"00",	-- Hex Addr	3523	13603
x"00",	-- Hex Addr	3524	13604
x"00",	-- Hex Addr	3525	13605
x"00",	-- Hex Addr	3526	13606
x"00",	-- Hex Addr	3527	13607
x"00",	-- Hex Addr	3528	13608
x"00",	-- Hex Addr	3529	13609
x"00",	-- Hex Addr	352A	13610
x"00",	-- Hex Addr	352B	13611
x"00",	-- Hex Addr	352C	13612
x"00",	-- Hex Addr	352D	13613
x"00",	-- Hex Addr	352E	13614
x"00",	-- Hex Addr	352F	13615
x"00",	-- Hex Addr	3530	13616
x"00",	-- Hex Addr	3531	13617
x"00",	-- Hex Addr	3532	13618
x"00",	-- Hex Addr	3533	13619
x"00",	-- Hex Addr	3534	13620
x"00",	-- Hex Addr	3535	13621
x"00",	-- Hex Addr	3536	13622
x"00",	-- Hex Addr	3537	13623
x"00",	-- Hex Addr	3538	13624
x"00",	-- Hex Addr	3539	13625
x"00",	-- Hex Addr	353A	13626
x"00",	-- Hex Addr	353B	13627
x"00",	-- Hex Addr	353C	13628
x"00",	-- Hex Addr	353D	13629
x"00",	-- Hex Addr	353E	13630
x"00",	-- Hex Addr	353F	13631
x"00",	-- Hex Addr	3540	13632
x"00",	-- Hex Addr	3541	13633
x"00",	-- Hex Addr	3542	13634
x"00",	-- Hex Addr	3543	13635
x"00",	-- Hex Addr	3544	13636
x"00",	-- Hex Addr	3545	13637
x"00",	-- Hex Addr	3546	13638
x"00",	-- Hex Addr	3547	13639
x"00",	-- Hex Addr	3548	13640
x"00",	-- Hex Addr	3549	13641
x"00",	-- Hex Addr	354A	13642
x"00",	-- Hex Addr	354B	13643
x"00",	-- Hex Addr	354C	13644
x"00",	-- Hex Addr	354D	13645
x"00",	-- Hex Addr	354E	13646
x"00",	-- Hex Addr	354F	13647
x"00",	-- Hex Addr	3550	13648
x"00",	-- Hex Addr	3551	13649
x"00",	-- Hex Addr	3552	13650
x"00",	-- Hex Addr	3553	13651
x"00",	-- Hex Addr	3554	13652
x"00",	-- Hex Addr	3555	13653
x"00",	-- Hex Addr	3556	13654
x"00",	-- Hex Addr	3557	13655
x"00",	-- Hex Addr	3558	13656
x"00",	-- Hex Addr	3559	13657
x"00",	-- Hex Addr	355A	13658
x"00",	-- Hex Addr	355B	13659
x"00",	-- Hex Addr	355C	13660
x"00",	-- Hex Addr	355D	13661
x"00",	-- Hex Addr	355E	13662
x"00",	-- Hex Addr	355F	13663
x"00",	-- Hex Addr	3560	13664
x"00",	-- Hex Addr	3561	13665
x"00",	-- Hex Addr	3562	13666
x"00",	-- Hex Addr	3563	13667
x"00",	-- Hex Addr	3564	13668
x"00",	-- Hex Addr	3565	13669
x"00",	-- Hex Addr	3566	13670
x"00",	-- Hex Addr	3567	13671
x"00",	-- Hex Addr	3568	13672
x"00",	-- Hex Addr	3569	13673
x"00",	-- Hex Addr	356A	13674
x"00",	-- Hex Addr	356B	13675
x"00",	-- Hex Addr	356C	13676
x"00",	-- Hex Addr	356D	13677
x"00",	-- Hex Addr	356E	13678
x"00",	-- Hex Addr	356F	13679
x"00",	-- Hex Addr	3570	13680
x"00",	-- Hex Addr	3571	13681
x"00",	-- Hex Addr	3572	13682
x"00",	-- Hex Addr	3573	13683
x"00",	-- Hex Addr	3574	13684
x"00",	-- Hex Addr	3575	13685
x"00",	-- Hex Addr	3576	13686
x"00",	-- Hex Addr	3577	13687
x"00",	-- Hex Addr	3578	13688
x"00",	-- Hex Addr	3579	13689
x"00",	-- Hex Addr	357A	13690
x"00",	-- Hex Addr	357B	13691
x"00",	-- Hex Addr	357C	13692
x"00",	-- Hex Addr	357D	13693
x"00",	-- Hex Addr	357E	13694
x"00",	-- Hex Addr	357F	13695
x"00",	-- Hex Addr	3580	13696
x"00",	-- Hex Addr	3581	13697
x"00",	-- Hex Addr	3582	13698
x"00",	-- Hex Addr	3583	13699
x"00",	-- Hex Addr	3584	13700
x"00",	-- Hex Addr	3585	13701
x"00",	-- Hex Addr	3586	13702
x"00",	-- Hex Addr	3587	13703
x"00",	-- Hex Addr	3588	13704
x"00",	-- Hex Addr	3589	13705
x"00",	-- Hex Addr	358A	13706
x"00",	-- Hex Addr	358B	13707
x"00",	-- Hex Addr	358C	13708
x"00",	-- Hex Addr	358D	13709
x"00",	-- Hex Addr	358E	13710
x"00",	-- Hex Addr	358F	13711
x"00",	-- Hex Addr	3590	13712
x"00",	-- Hex Addr	3591	13713
x"00",	-- Hex Addr	3592	13714
x"00",	-- Hex Addr	3593	13715
x"00",	-- Hex Addr	3594	13716
x"00",	-- Hex Addr	3595	13717
x"00",	-- Hex Addr	3596	13718
x"00",	-- Hex Addr	3597	13719
x"00",	-- Hex Addr	3598	13720
x"00",	-- Hex Addr	3599	13721
x"00",	-- Hex Addr	359A	13722
x"00",	-- Hex Addr	359B	13723
x"00",	-- Hex Addr	359C	13724
x"00",	-- Hex Addr	359D	13725
x"00",	-- Hex Addr	359E	13726
x"00",	-- Hex Addr	359F	13727
x"00",	-- Hex Addr	35A0	13728
x"00",	-- Hex Addr	35A1	13729
x"00",	-- Hex Addr	35A2	13730
x"00",	-- Hex Addr	35A3	13731
x"00",	-- Hex Addr	35A4	13732
x"00",	-- Hex Addr	35A5	13733
x"00",	-- Hex Addr	35A6	13734
x"00",	-- Hex Addr	35A7	13735
x"00",	-- Hex Addr	35A8	13736
x"00",	-- Hex Addr	35A9	13737
x"00",	-- Hex Addr	35AA	13738
x"00",	-- Hex Addr	35AB	13739
x"00",	-- Hex Addr	35AC	13740
x"00",	-- Hex Addr	35AD	13741
x"00",	-- Hex Addr	35AE	13742
x"00",	-- Hex Addr	35AF	13743
x"00",	-- Hex Addr	35B0	13744
x"00",	-- Hex Addr	35B1	13745
x"00",	-- Hex Addr	35B2	13746
x"00",	-- Hex Addr	35B3	13747
x"00",	-- Hex Addr	35B4	13748
x"00",	-- Hex Addr	35B5	13749
x"00",	-- Hex Addr	35B6	13750
x"00",	-- Hex Addr	35B7	13751
x"00",	-- Hex Addr	35B8	13752
x"00",	-- Hex Addr	35B9	13753
x"00",	-- Hex Addr	35BA	13754
x"00",	-- Hex Addr	35BB	13755
x"00",	-- Hex Addr	35BC	13756
x"00",	-- Hex Addr	35BD	13757
x"00",	-- Hex Addr	35BE	13758
x"00",	-- Hex Addr	35BF	13759
x"00",	-- Hex Addr	35C0	13760
x"00",	-- Hex Addr	35C1	13761
x"00",	-- Hex Addr	35C2	13762
x"00",	-- Hex Addr	35C3	13763
x"00",	-- Hex Addr	35C4	13764
x"00",	-- Hex Addr	35C5	13765
x"00",	-- Hex Addr	35C6	13766
x"00",	-- Hex Addr	35C7	13767
x"00",	-- Hex Addr	35C8	13768
x"00",	-- Hex Addr	35C9	13769
x"00",	-- Hex Addr	35CA	13770
x"00",	-- Hex Addr	35CB	13771
x"00",	-- Hex Addr	35CC	13772
x"00",	-- Hex Addr	35CD	13773
x"00",	-- Hex Addr	35CE	13774
x"00",	-- Hex Addr	35CF	13775
x"00",	-- Hex Addr	35D0	13776
x"00",	-- Hex Addr	35D1	13777
x"00",	-- Hex Addr	35D2	13778
x"00",	-- Hex Addr	35D3	13779
x"00",	-- Hex Addr	35D4	13780
x"00",	-- Hex Addr	35D5	13781
x"00",	-- Hex Addr	35D6	13782
x"00",	-- Hex Addr	35D7	13783
x"00",	-- Hex Addr	35D8	13784
x"00",	-- Hex Addr	35D9	13785
x"00",	-- Hex Addr	35DA	13786
x"00",	-- Hex Addr	35DB	13787
x"00",	-- Hex Addr	35DC	13788
x"00",	-- Hex Addr	35DD	13789
x"00",	-- Hex Addr	35DE	13790
x"00",	-- Hex Addr	35DF	13791
x"00",	-- Hex Addr	35E0	13792
x"00",	-- Hex Addr	35E1	13793
x"00",	-- Hex Addr	35E2	13794
x"00",	-- Hex Addr	35E3	13795
x"00",	-- Hex Addr	35E4	13796
x"00",	-- Hex Addr	35E5	13797
x"00",	-- Hex Addr	35E6	13798
x"00",	-- Hex Addr	35E7	13799
x"00",	-- Hex Addr	35E8	13800
x"00",	-- Hex Addr	35E9	13801
x"00",	-- Hex Addr	35EA	13802
x"00",	-- Hex Addr	35EB	13803
x"00",	-- Hex Addr	35EC	13804
x"00",	-- Hex Addr	35ED	13805
x"00",	-- Hex Addr	35EE	13806
x"00",	-- Hex Addr	35EF	13807
x"00",	-- Hex Addr	35F0	13808
x"00",	-- Hex Addr	35F1	13809
x"00",	-- Hex Addr	35F2	13810
x"00",	-- Hex Addr	35F3	13811
x"00",	-- Hex Addr	35F4	13812
x"00",	-- Hex Addr	35F5	13813
x"00",	-- Hex Addr	35F6	13814
x"00",	-- Hex Addr	35F7	13815
x"00",	-- Hex Addr	35F8	13816
x"00",	-- Hex Addr	35F9	13817
x"00",	-- Hex Addr	35FA	13818
x"00",	-- Hex Addr	35FB	13819
x"00",	-- Hex Addr	35FC	13820
x"00",	-- Hex Addr	35FD	13821
x"00",	-- Hex Addr	35FE	13822
x"00",	-- Hex Addr	35FF	13823
x"00",	-- Hex Addr	3600	13824
x"00",	-- Hex Addr	3601	13825
x"00",	-- Hex Addr	3602	13826
x"00",	-- Hex Addr	3603	13827
x"00",	-- Hex Addr	3604	13828
x"00",	-- Hex Addr	3605	13829
x"00",	-- Hex Addr	3606	13830
x"00",	-- Hex Addr	3607	13831
x"00",	-- Hex Addr	3608	13832
x"00",	-- Hex Addr	3609	13833
x"00",	-- Hex Addr	360A	13834
x"00",	-- Hex Addr	360B	13835
x"00",	-- Hex Addr	360C	13836
x"00",	-- Hex Addr	360D	13837
x"00",	-- Hex Addr	360E	13838
x"00",	-- Hex Addr	360F	13839
x"00",	-- Hex Addr	3610	13840
x"00",	-- Hex Addr	3611	13841
x"00",	-- Hex Addr	3612	13842
x"00",	-- Hex Addr	3613	13843
x"00",	-- Hex Addr	3614	13844
x"00",	-- Hex Addr	3615	13845
x"00",	-- Hex Addr	3616	13846
x"00",	-- Hex Addr	3617	13847
x"00",	-- Hex Addr	3618	13848
x"00",	-- Hex Addr	3619	13849
x"00",	-- Hex Addr	361A	13850
x"00",	-- Hex Addr	361B	13851
x"00",	-- Hex Addr	361C	13852
x"00",	-- Hex Addr	361D	13853
x"00",	-- Hex Addr	361E	13854
x"00",	-- Hex Addr	361F	13855
x"00",	-- Hex Addr	3620	13856
x"00",	-- Hex Addr	3621	13857
x"00",	-- Hex Addr	3622	13858
x"00",	-- Hex Addr	3623	13859
x"00",	-- Hex Addr	3624	13860
x"00",	-- Hex Addr	3625	13861
x"00",	-- Hex Addr	3626	13862
x"00",	-- Hex Addr	3627	13863
x"00",	-- Hex Addr	3628	13864
x"00",	-- Hex Addr	3629	13865
x"00",	-- Hex Addr	362A	13866
x"00",	-- Hex Addr	362B	13867
x"00",	-- Hex Addr	362C	13868
x"00",	-- Hex Addr	362D	13869
x"00",	-- Hex Addr	362E	13870
x"00",	-- Hex Addr	362F	13871
x"00",	-- Hex Addr	3630	13872
x"00",	-- Hex Addr	3631	13873
x"00",	-- Hex Addr	3632	13874
x"00",	-- Hex Addr	3633	13875
x"00",	-- Hex Addr	3634	13876
x"00",	-- Hex Addr	3635	13877
x"00",	-- Hex Addr	3636	13878
x"00",	-- Hex Addr	3637	13879
x"00",	-- Hex Addr	3638	13880
x"00",	-- Hex Addr	3639	13881
x"00",	-- Hex Addr	363A	13882
x"00",	-- Hex Addr	363B	13883
x"00",	-- Hex Addr	363C	13884
x"00",	-- Hex Addr	363D	13885
x"00",	-- Hex Addr	363E	13886
x"00",	-- Hex Addr	363F	13887
x"00",	-- Hex Addr	3640	13888
x"00",	-- Hex Addr	3641	13889
x"00",	-- Hex Addr	3642	13890
x"00",	-- Hex Addr	3643	13891
x"00",	-- Hex Addr	3644	13892
x"00",	-- Hex Addr	3645	13893
x"00",	-- Hex Addr	3646	13894
x"00",	-- Hex Addr	3647	13895
x"00",	-- Hex Addr	3648	13896
x"00",	-- Hex Addr	3649	13897
x"00",	-- Hex Addr	364A	13898
x"00",	-- Hex Addr	364B	13899
x"00",	-- Hex Addr	364C	13900
x"00",	-- Hex Addr	364D	13901
x"00",	-- Hex Addr	364E	13902
x"00",	-- Hex Addr	364F	13903
x"00",	-- Hex Addr	3650	13904
x"00",	-- Hex Addr	3651	13905
x"00",	-- Hex Addr	3652	13906
x"00",	-- Hex Addr	3653	13907
x"00",	-- Hex Addr	3654	13908
x"00",	-- Hex Addr	3655	13909
x"00",	-- Hex Addr	3656	13910
x"00",	-- Hex Addr	3657	13911
x"00",	-- Hex Addr	3658	13912
x"00",	-- Hex Addr	3659	13913
x"00",	-- Hex Addr	365A	13914
x"00",	-- Hex Addr	365B	13915
x"00",	-- Hex Addr	365C	13916
x"00",	-- Hex Addr	365D	13917
x"00",	-- Hex Addr	365E	13918
x"00",	-- Hex Addr	365F	13919
x"00",	-- Hex Addr	3660	13920
x"00",	-- Hex Addr	3661	13921
x"00",	-- Hex Addr	3662	13922
x"00",	-- Hex Addr	3663	13923
x"00",	-- Hex Addr	3664	13924
x"00",	-- Hex Addr	3665	13925
x"00",	-- Hex Addr	3666	13926
x"00",	-- Hex Addr	3667	13927
x"00",	-- Hex Addr	3668	13928
x"00",	-- Hex Addr	3669	13929
x"00",	-- Hex Addr	366A	13930
x"00",	-- Hex Addr	366B	13931
x"00",	-- Hex Addr	366C	13932
x"00",	-- Hex Addr	366D	13933
x"00",	-- Hex Addr	366E	13934
x"00",	-- Hex Addr	366F	13935
x"00",	-- Hex Addr	3670	13936
x"00",	-- Hex Addr	3671	13937
x"00",	-- Hex Addr	3672	13938
x"00",	-- Hex Addr	3673	13939
x"00",	-- Hex Addr	3674	13940
x"00",	-- Hex Addr	3675	13941
x"00",	-- Hex Addr	3676	13942
x"00",	-- Hex Addr	3677	13943
x"00",	-- Hex Addr	3678	13944
x"00",	-- Hex Addr	3679	13945
x"00",	-- Hex Addr	367A	13946
x"00",	-- Hex Addr	367B	13947
x"00",	-- Hex Addr	367C	13948
x"00",	-- Hex Addr	367D	13949
x"00",	-- Hex Addr	367E	13950
x"00",	-- Hex Addr	367F	13951
x"00",	-- Hex Addr	3680	13952
x"00",	-- Hex Addr	3681	13953
x"00",	-- Hex Addr	3682	13954
x"00",	-- Hex Addr	3683	13955
x"00",	-- Hex Addr	3684	13956
x"00",	-- Hex Addr	3685	13957
x"00",	-- Hex Addr	3686	13958
x"00",	-- Hex Addr	3687	13959
x"00",	-- Hex Addr	3688	13960
x"00",	-- Hex Addr	3689	13961
x"00",	-- Hex Addr	368A	13962
x"00",	-- Hex Addr	368B	13963
x"00",	-- Hex Addr	368C	13964
x"00",	-- Hex Addr	368D	13965
x"00",	-- Hex Addr	368E	13966
x"00",	-- Hex Addr	368F	13967
x"00",	-- Hex Addr	3690	13968
x"00",	-- Hex Addr	3691	13969
x"00",	-- Hex Addr	3692	13970
x"00",	-- Hex Addr	3693	13971
x"00",	-- Hex Addr	3694	13972
x"00",	-- Hex Addr	3695	13973
x"00",	-- Hex Addr	3696	13974
x"00",	-- Hex Addr	3697	13975
x"00",	-- Hex Addr	3698	13976
x"00",	-- Hex Addr	3699	13977
x"00",	-- Hex Addr	369A	13978
x"00",	-- Hex Addr	369B	13979
x"00",	-- Hex Addr	369C	13980
x"00",	-- Hex Addr	369D	13981
x"00",	-- Hex Addr	369E	13982
x"00",	-- Hex Addr	369F	13983
x"00",	-- Hex Addr	36A0	13984
x"00",	-- Hex Addr	36A1	13985
x"00",	-- Hex Addr	36A2	13986
x"00",	-- Hex Addr	36A3	13987
x"00",	-- Hex Addr	36A4	13988
x"00",	-- Hex Addr	36A5	13989
x"00",	-- Hex Addr	36A6	13990
x"00",	-- Hex Addr	36A7	13991
x"00",	-- Hex Addr	36A8	13992
x"00",	-- Hex Addr	36A9	13993
x"00",	-- Hex Addr	36AA	13994
x"00",	-- Hex Addr	36AB	13995
x"00",	-- Hex Addr	36AC	13996
x"00",	-- Hex Addr	36AD	13997
x"00",	-- Hex Addr	36AE	13998
x"00",	-- Hex Addr	36AF	13999
x"00",	-- Hex Addr	36B0	14000
x"00",	-- Hex Addr	36B1	14001
x"00",	-- Hex Addr	36B2	14002
x"00",	-- Hex Addr	36B3	14003
x"00",	-- Hex Addr	36B4	14004
x"00",	-- Hex Addr	36B5	14005
x"00",	-- Hex Addr	36B6	14006
x"00",	-- Hex Addr	36B7	14007
x"00",	-- Hex Addr	36B8	14008
x"00",	-- Hex Addr	36B9	14009
x"00",	-- Hex Addr	36BA	14010
x"00",	-- Hex Addr	36BB	14011
x"00",	-- Hex Addr	36BC	14012
x"00",	-- Hex Addr	36BD	14013
x"00",	-- Hex Addr	36BE	14014
x"00",	-- Hex Addr	36BF	14015
x"00",	-- Hex Addr	36C0	14016
x"00",	-- Hex Addr	36C1	14017
x"00",	-- Hex Addr	36C2	14018
x"00",	-- Hex Addr	36C3	14019
x"00",	-- Hex Addr	36C4	14020
x"00",	-- Hex Addr	36C5	14021
x"00",	-- Hex Addr	36C6	14022
x"00",	-- Hex Addr	36C7	14023
x"00",	-- Hex Addr	36C8	14024
x"00",	-- Hex Addr	36C9	14025
x"00",	-- Hex Addr	36CA	14026
x"00",	-- Hex Addr	36CB	14027
x"00",	-- Hex Addr	36CC	14028
x"00",	-- Hex Addr	36CD	14029
x"00",	-- Hex Addr	36CE	14030
x"00",	-- Hex Addr	36CF	14031
x"00",	-- Hex Addr	36D0	14032
x"00",	-- Hex Addr	36D1	14033
x"00",	-- Hex Addr	36D2	14034
x"00",	-- Hex Addr	36D3	14035
x"00",	-- Hex Addr	36D4	14036
x"00",	-- Hex Addr	36D5	14037
x"00",	-- Hex Addr	36D6	14038
x"00",	-- Hex Addr	36D7	14039
x"00",	-- Hex Addr	36D8	14040
x"00",	-- Hex Addr	36D9	14041
x"00",	-- Hex Addr	36DA	14042
x"00",	-- Hex Addr	36DB	14043
x"00",	-- Hex Addr	36DC	14044
x"00",	-- Hex Addr	36DD	14045
x"00",	-- Hex Addr	36DE	14046
x"00",	-- Hex Addr	36DF	14047
x"00",	-- Hex Addr	36E0	14048
x"00",	-- Hex Addr	36E1	14049
x"00",	-- Hex Addr	36E2	14050
x"00",	-- Hex Addr	36E3	14051
x"00",	-- Hex Addr	36E4	14052
x"00",	-- Hex Addr	36E5	14053
x"00",	-- Hex Addr	36E6	14054
x"00",	-- Hex Addr	36E7	14055
x"00",	-- Hex Addr	36E8	14056
x"00",	-- Hex Addr	36E9	14057
x"00",	-- Hex Addr	36EA	14058
x"00",	-- Hex Addr	36EB	14059
x"00",	-- Hex Addr	36EC	14060
x"00",	-- Hex Addr	36ED	14061
x"00",	-- Hex Addr	36EE	14062
x"00",	-- Hex Addr	36EF	14063
x"00",	-- Hex Addr	36F0	14064
x"00",	-- Hex Addr	36F1	14065
x"00",	-- Hex Addr	36F2	14066
x"00",	-- Hex Addr	36F3	14067
x"00",	-- Hex Addr	36F4	14068
x"00",	-- Hex Addr	36F5	14069
x"00",	-- Hex Addr	36F6	14070
x"00",	-- Hex Addr	36F7	14071
x"00",	-- Hex Addr	36F8	14072
x"00",	-- Hex Addr	36F9	14073
x"00",	-- Hex Addr	36FA	14074
x"00",	-- Hex Addr	36FB	14075
x"00",	-- Hex Addr	36FC	14076
x"00",	-- Hex Addr	36FD	14077
x"00",	-- Hex Addr	36FE	14078
x"00",	-- Hex Addr	36FF	14079
x"00",	-- Hex Addr	3700	14080
x"00",	-- Hex Addr	3701	14081
x"00",	-- Hex Addr	3702	14082
x"00",	-- Hex Addr	3703	14083
x"00",	-- Hex Addr	3704	14084
x"00",	-- Hex Addr	3705	14085
x"00",	-- Hex Addr	3706	14086
x"00",	-- Hex Addr	3707	14087
x"00",	-- Hex Addr	3708	14088
x"00",	-- Hex Addr	3709	14089
x"00",	-- Hex Addr	370A	14090
x"00",	-- Hex Addr	370B	14091
x"00",	-- Hex Addr	370C	14092
x"00",	-- Hex Addr	370D	14093
x"00",	-- Hex Addr	370E	14094
x"00",	-- Hex Addr	370F	14095
x"00",	-- Hex Addr	3710	14096
x"00",	-- Hex Addr	3711	14097
x"00",	-- Hex Addr	3712	14098
x"00",	-- Hex Addr	3713	14099
x"00",	-- Hex Addr	3714	14100
x"00",	-- Hex Addr	3715	14101
x"00",	-- Hex Addr	3716	14102
x"00",	-- Hex Addr	3717	14103
x"00",	-- Hex Addr	3718	14104
x"00",	-- Hex Addr	3719	14105
x"00",	-- Hex Addr	371A	14106
x"00",	-- Hex Addr	371B	14107
x"00",	-- Hex Addr	371C	14108
x"00",	-- Hex Addr	371D	14109
x"00",	-- Hex Addr	371E	14110
x"00",	-- Hex Addr	371F	14111
x"00",	-- Hex Addr	3720	14112
x"00",	-- Hex Addr	3721	14113
x"00",	-- Hex Addr	3722	14114
x"00",	-- Hex Addr	3723	14115
x"00",	-- Hex Addr	3724	14116
x"00",	-- Hex Addr	3725	14117
x"00",	-- Hex Addr	3726	14118
x"00",	-- Hex Addr	3727	14119
x"00",	-- Hex Addr	3728	14120
x"00",	-- Hex Addr	3729	14121
x"00",	-- Hex Addr	372A	14122
x"00",	-- Hex Addr	372B	14123
x"00",	-- Hex Addr	372C	14124
x"00",	-- Hex Addr	372D	14125
x"00",	-- Hex Addr	372E	14126
x"00",	-- Hex Addr	372F	14127
x"00",	-- Hex Addr	3730	14128
x"00",	-- Hex Addr	3731	14129
x"00",	-- Hex Addr	3732	14130
x"00",	-- Hex Addr	3733	14131
x"00",	-- Hex Addr	3734	14132
x"00",	-- Hex Addr	3735	14133
x"00",	-- Hex Addr	3736	14134
x"00",	-- Hex Addr	3737	14135
x"00",	-- Hex Addr	3738	14136
x"00",	-- Hex Addr	3739	14137
x"00",	-- Hex Addr	373A	14138
x"00",	-- Hex Addr	373B	14139
x"00",	-- Hex Addr	373C	14140
x"00",	-- Hex Addr	373D	14141
x"00",	-- Hex Addr	373E	14142
x"00",	-- Hex Addr	373F	14143
x"00",	-- Hex Addr	3740	14144
x"00",	-- Hex Addr	3741	14145
x"00",	-- Hex Addr	3742	14146
x"00",	-- Hex Addr	3743	14147
x"00",	-- Hex Addr	3744	14148
x"00",	-- Hex Addr	3745	14149
x"00",	-- Hex Addr	3746	14150
x"00",	-- Hex Addr	3747	14151
x"00",	-- Hex Addr	3748	14152
x"00",	-- Hex Addr	3749	14153
x"00",	-- Hex Addr	374A	14154
x"00",	-- Hex Addr	374B	14155
x"00",	-- Hex Addr	374C	14156
x"00",	-- Hex Addr	374D	14157
x"00",	-- Hex Addr	374E	14158
x"00",	-- Hex Addr	374F	14159
x"00",	-- Hex Addr	3750	14160
x"00",	-- Hex Addr	3751	14161
x"00",	-- Hex Addr	3752	14162
x"00",	-- Hex Addr	3753	14163
x"00",	-- Hex Addr	3754	14164
x"00",	-- Hex Addr	3755	14165
x"00",	-- Hex Addr	3756	14166
x"00",	-- Hex Addr	3757	14167
x"00",	-- Hex Addr	3758	14168
x"00",	-- Hex Addr	3759	14169
x"00",	-- Hex Addr	375A	14170
x"00",	-- Hex Addr	375B	14171
x"00",	-- Hex Addr	375C	14172
x"00",	-- Hex Addr	375D	14173
x"00",	-- Hex Addr	375E	14174
x"00",	-- Hex Addr	375F	14175
x"00",	-- Hex Addr	3760	14176
x"00",	-- Hex Addr	3761	14177
x"00",	-- Hex Addr	3762	14178
x"00",	-- Hex Addr	3763	14179
x"00",	-- Hex Addr	3764	14180
x"00",	-- Hex Addr	3765	14181
x"00",	-- Hex Addr	3766	14182
x"00",	-- Hex Addr	3767	14183
x"00",	-- Hex Addr	3768	14184
x"00",	-- Hex Addr	3769	14185
x"00",	-- Hex Addr	376A	14186
x"00",	-- Hex Addr	376B	14187
x"00",	-- Hex Addr	376C	14188
x"00",	-- Hex Addr	376D	14189
x"00",	-- Hex Addr	376E	14190
x"00",	-- Hex Addr	376F	14191
x"00",	-- Hex Addr	3770	14192
x"00",	-- Hex Addr	3771	14193
x"00",	-- Hex Addr	3772	14194
x"00",	-- Hex Addr	3773	14195
x"00",	-- Hex Addr	3774	14196
x"00",	-- Hex Addr	3775	14197
x"00",	-- Hex Addr	3776	14198
x"00",	-- Hex Addr	3777	14199
x"00",	-- Hex Addr	3778	14200
x"00",	-- Hex Addr	3779	14201
x"00",	-- Hex Addr	377A	14202
x"00",	-- Hex Addr	377B	14203
x"00",	-- Hex Addr	377C	14204
x"00",	-- Hex Addr	377D	14205
x"00",	-- Hex Addr	377E	14206
x"00",	-- Hex Addr	377F	14207
x"00",	-- Hex Addr	3780	14208
x"00",	-- Hex Addr	3781	14209
x"00",	-- Hex Addr	3782	14210
x"00",	-- Hex Addr	3783	14211
x"00",	-- Hex Addr	3784	14212
x"00",	-- Hex Addr	3785	14213
x"00",	-- Hex Addr	3786	14214
x"00",	-- Hex Addr	3787	14215
x"00",	-- Hex Addr	3788	14216
x"00",	-- Hex Addr	3789	14217
x"00",	-- Hex Addr	378A	14218
x"00",	-- Hex Addr	378B	14219
x"00",	-- Hex Addr	378C	14220
x"00",	-- Hex Addr	378D	14221
x"00",	-- Hex Addr	378E	14222
x"00",	-- Hex Addr	378F	14223
x"00",	-- Hex Addr	3790	14224
x"00",	-- Hex Addr	3791	14225
x"00",	-- Hex Addr	3792	14226
x"00",	-- Hex Addr	3793	14227
x"00",	-- Hex Addr	3794	14228
x"00",	-- Hex Addr	3795	14229
x"00",	-- Hex Addr	3796	14230
x"00",	-- Hex Addr	3797	14231
x"00",	-- Hex Addr	3798	14232
x"00",	-- Hex Addr	3799	14233
x"00",	-- Hex Addr	379A	14234
x"00",	-- Hex Addr	379B	14235
x"00",	-- Hex Addr	379C	14236
x"00",	-- Hex Addr	379D	14237
x"00",	-- Hex Addr	379E	14238
x"00",	-- Hex Addr	379F	14239
x"00",	-- Hex Addr	37A0	14240
x"00",	-- Hex Addr	37A1	14241
x"00",	-- Hex Addr	37A2	14242
x"00",	-- Hex Addr	37A3	14243
x"00",	-- Hex Addr	37A4	14244
x"00",	-- Hex Addr	37A5	14245
x"00",	-- Hex Addr	37A6	14246
x"00",	-- Hex Addr	37A7	14247
x"00",	-- Hex Addr	37A8	14248
x"00",	-- Hex Addr	37A9	14249
x"00",	-- Hex Addr	37AA	14250
x"00",	-- Hex Addr	37AB	14251
x"00",	-- Hex Addr	37AC	14252
x"00",	-- Hex Addr	37AD	14253
x"00",	-- Hex Addr	37AE	14254
x"00",	-- Hex Addr	37AF	14255
x"00",	-- Hex Addr	37B0	14256
x"00",	-- Hex Addr	37B1	14257
x"00",	-- Hex Addr	37B2	14258
x"00",	-- Hex Addr	37B3	14259
x"00",	-- Hex Addr	37B4	14260
x"00",	-- Hex Addr	37B5	14261
x"00",	-- Hex Addr	37B6	14262
x"00",	-- Hex Addr	37B7	14263
x"00",	-- Hex Addr	37B8	14264
x"00",	-- Hex Addr	37B9	14265
x"00",	-- Hex Addr	37BA	14266
x"00",	-- Hex Addr	37BB	14267
x"00",	-- Hex Addr	37BC	14268
x"00",	-- Hex Addr	37BD	14269
x"00",	-- Hex Addr	37BE	14270
x"00",	-- Hex Addr	37BF	14271
x"00",	-- Hex Addr	37C0	14272
x"00",	-- Hex Addr	37C1	14273
x"00",	-- Hex Addr	37C2	14274
x"00",	-- Hex Addr	37C3	14275
x"00",	-- Hex Addr	37C4	14276
x"00",	-- Hex Addr	37C5	14277
x"00",	-- Hex Addr	37C6	14278
x"00",	-- Hex Addr	37C7	14279
x"00",	-- Hex Addr	37C8	14280
x"00",	-- Hex Addr	37C9	14281
x"00",	-- Hex Addr	37CA	14282
x"00",	-- Hex Addr	37CB	14283
x"00",	-- Hex Addr	37CC	14284
x"00",	-- Hex Addr	37CD	14285
x"00",	-- Hex Addr	37CE	14286
x"00",	-- Hex Addr	37CF	14287
x"00",	-- Hex Addr	37D0	14288
x"00",	-- Hex Addr	37D1	14289
x"00",	-- Hex Addr	37D2	14290
x"00",	-- Hex Addr	37D3	14291
x"00",	-- Hex Addr	37D4	14292
x"00",	-- Hex Addr	37D5	14293
x"00",	-- Hex Addr	37D6	14294
x"00",	-- Hex Addr	37D7	14295
x"00",	-- Hex Addr	37D8	14296
x"00",	-- Hex Addr	37D9	14297
x"00",	-- Hex Addr	37DA	14298
x"00",	-- Hex Addr	37DB	14299
x"00",	-- Hex Addr	37DC	14300
x"00",	-- Hex Addr	37DD	14301
x"00",	-- Hex Addr	37DE	14302
x"00",	-- Hex Addr	37DF	14303
x"00",	-- Hex Addr	37E0	14304
x"00",	-- Hex Addr	37E1	14305
x"00",	-- Hex Addr	37E2	14306
x"00",	-- Hex Addr	37E3	14307
x"00",	-- Hex Addr	37E4	14308
x"00",	-- Hex Addr	37E5	14309
x"00",	-- Hex Addr	37E6	14310
x"00",	-- Hex Addr	37E7	14311
x"00",	-- Hex Addr	37E8	14312
x"00",	-- Hex Addr	37E9	14313
x"00",	-- Hex Addr	37EA	14314
x"00",	-- Hex Addr	37EB	14315
x"00",	-- Hex Addr	37EC	14316
x"00",	-- Hex Addr	37ED	14317
x"00",	-- Hex Addr	37EE	14318
x"00",	-- Hex Addr	37EF	14319
x"00",	-- Hex Addr	37F0	14320
x"00",	-- Hex Addr	37F1	14321
x"00",	-- Hex Addr	37F2	14322
x"00",	-- Hex Addr	37F3	14323
x"00",	-- Hex Addr	37F4	14324
x"00",	-- Hex Addr	37F5	14325
x"00",	-- Hex Addr	37F6	14326
x"00",	-- Hex Addr	37F7	14327
x"00",	-- Hex Addr	37F8	14328
x"00",	-- Hex Addr	37F9	14329
x"00",	-- Hex Addr	37FA	14330
x"00",	-- Hex Addr	37FB	14331
x"00",	-- Hex Addr	37FC	14332
x"00",	-- Hex Addr	37FD	14333
x"00",	-- Hex Addr	37FE	14334
x"00",	-- Hex Addr	37FF	14335
x"00",	-- Hex Addr	3800	14336
x"00",	-- Hex Addr	3801	14337
x"00",	-- Hex Addr	3802	14338
x"00",	-- Hex Addr	3803	14339
x"00",	-- Hex Addr	3804	14340
x"00",	-- Hex Addr	3805	14341
x"00",	-- Hex Addr	3806	14342
x"00",	-- Hex Addr	3807	14343
x"00",	-- Hex Addr	3808	14344
x"00",	-- Hex Addr	3809	14345
x"00",	-- Hex Addr	380A	14346
x"00",	-- Hex Addr	380B	14347
x"00",	-- Hex Addr	380C	14348
x"00",	-- Hex Addr	380D	14349
x"00",	-- Hex Addr	380E	14350
x"00",	-- Hex Addr	380F	14351
x"00",	-- Hex Addr	3810	14352
x"00",	-- Hex Addr	3811	14353
x"00",	-- Hex Addr	3812	14354
x"00",	-- Hex Addr	3813	14355
x"00",	-- Hex Addr	3814	14356
x"00",	-- Hex Addr	3815	14357
x"00",	-- Hex Addr	3816	14358
x"00",	-- Hex Addr	3817	14359
x"00",	-- Hex Addr	3818	14360
x"00",	-- Hex Addr	3819	14361
x"00",	-- Hex Addr	381A	14362
x"00",	-- Hex Addr	381B	14363
x"00",	-- Hex Addr	381C	14364
x"00",	-- Hex Addr	381D	14365
x"00",	-- Hex Addr	381E	14366
x"00",	-- Hex Addr	381F	14367
x"00",	-- Hex Addr	3820	14368
x"00",	-- Hex Addr	3821	14369
x"00",	-- Hex Addr	3822	14370
x"00",	-- Hex Addr	3823	14371
x"00",	-- Hex Addr	3824	14372
x"00",	-- Hex Addr	3825	14373
x"00",	-- Hex Addr	3826	14374
x"00",	-- Hex Addr	3827	14375
x"00",	-- Hex Addr	3828	14376
x"00",	-- Hex Addr	3829	14377
x"00",	-- Hex Addr	382A	14378
x"00",	-- Hex Addr	382B	14379
x"00",	-- Hex Addr	382C	14380
x"00",	-- Hex Addr	382D	14381
x"00",	-- Hex Addr	382E	14382
x"00",	-- Hex Addr	382F	14383
x"00",	-- Hex Addr	3830	14384
x"00",	-- Hex Addr	3831	14385
x"00",	-- Hex Addr	3832	14386
x"00",	-- Hex Addr	3833	14387
x"00",	-- Hex Addr	3834	14388
x"00",	-- Hex Addr	3835	14389
x"00",	-- Hex Addr	3836	14390
x"00",	-- Hex Addr	3837	14391
x"00",	-- Hex Addr	3838	14392
x"00",	-- Hex Addr	3839	14393
x"00",	-- Hex Addr	383A	14394
x"00",	-- Hex Addr	383B	14395
x"00",	-- Hex Addr	383C	14396
x"00",	-- Hex Addr	383D	14397
x"00",	-- Hex Addr	383E	14398
x"00",	-- Hex Addr	383F	14399
x"00",	-- Hex Addr	3840	14400
x"00",	-- Hex Addr	3841	14401
x"00",	-- Hex Addr	3842	14402
x"00",	-- Hex Addr	3843	14403
x"00",	-- Hex Addr	3844	14404
x"00",	-- Hex Addr	3845	14405
x"00",	-- Hex Addr	3846	14406
x"00",	-- Hex Addr	3847	14407
x"00",	-- Hex Addr	3848	14408
x"00",	-- Hex Addr	3849	14409
x"00",	-- Hex Addr	384A	14410
x"00",	-- Hex Addr	384B	14411
x"00",	-- Hex Addr	384C	14412
x"00",	-- Hex Addr	384D	14413
x"00",	-- Hex Addr	384E	14414
x"00",	-- Hex Addr	384F	14415
x"00",	-- Hex Addr	3850	14416
x"00",	-- Hex Addr	3851	14417
x"00",	-- Hex Addr	3852	14418
x"00",	-- Hex Addr	3853	14419
x"00",	-- Hex Addr	3854	14420
x"00",	-- Hex Addr	3855	14421
x"00",	-- Hex Addr	3856	14422
x"00",	-- Hex Addr	3857	14423
x"00",	-- Hex Addr	3858	14424
x"00",	-- Hex Addr	3859	14425
x"00",	-- Hex Addr	385A	14426
x"00",	-- Hex Addr	385B	14427
x"00",	-- Hex Addr	385C	14428
x"00",	-- Hex Addr	385D	14429
x"00",	-- Hex Addr	385E	14430
x"00",	-- Hex Addr	385F	14431
x"00",	-- Hex Addr	3860	14432
x"00",	-- Hex Addr	3861	14433
x"00",	-- Hex Addr	3862	14434
x"00",	-- Hex Addr	3863	14435
x"00",	-- Hex Addr	3864	14436
x"00",	-- Hex Addr	3865	14437
x"00",	-- Hex Addr	3866	14438
x"00",	-- Hex Addr	3867	14439
x"00",	-- Hex Addr	3868	14440
x"00",	-- Hex Addr	3869	14441
x"00",	-- Hex Addr	386A	14442
x"00",	-- Hex Addr	386B	14443
x"00",	-- Hex Addr	386C	14444
x"00",	-- Hex Addr	386D	14445
x"00",	-- Hex Addr	386E	14446
x"00",	-- Hex Addr	386F	14447
x"00",	-- Hex Addr	3870	14448
x"00",	-- Hex Addr	3871	14449
x"00",	-- Hex Addr	3872	14450
x"00",	-- Hex Addr	3873	14451
x"00",	-- Hex Addr	3874	14452
x"00",	-- Hex Addr	3875	14453
x"00",	-- Hex Addr	3876	14454
x"00",	-- Hex Addr	3877	14455
x"00",	-- Hex Addr	3878	14456
x"00",	-- Hex Addr	3879	14457
x"00",	-- Hex Addr	387A	14458
x"00",	-- Hex Addr	387B	14459
x"00",	-- Hex Addr	387C	14460
x"00",	-- Hex Addr	387D	14461
x"00",	-- Hex Addr	387E	14462
x"00",	-- Hex Addr	387F	14463
x"00",	-- Hex Addr	3880	14464
x"00",	-- Hex Addr	3881	14465
x"00",	-- Hex Addr	3882	14466
x"00",	-- Hex Addr	3883	14467
x"00",	-- Hex Addr	3884	14468
x"00",	-- Hex Addr	3885	14469
x"00",	-- Hex Addr	3886	14470
x"00",	-- Hex Addr	3887	14471
x"00",	-- Hex Addr	3888	14472
x"00",	-- Hex Addr	3889	14473
x"00",	-- Hex Addr	388A	14474
x"00",	-- Hex Addr	388B	14475
x"00",	-- Hex Addr	388C	14476
x"00",	-- Hex Addr	388D	14477
x"00",	-- Hex Addr	388E	14478
x"00",	-- Hex Addr	388F	14479
x"00",	-- Hex Addr	3890	14480
x"00",	-- Hex Addr	3891	14481
x"00",	-- Hex Addr	3892	14482
x"00",	-- Hex Addr	3893	14483
x"00",	-- Hex Addr	3894	14484
x"00",	-- Hex Addr	3895	14485
x"00",	-- Hex Addr	3896	14486
x"00",	-- Hex Addr	3897	14487
x"00",	-- Hex Addr	3898	14488
x"00",	-- Hex Addr	3899	14489
x"00",	-- Hex Addr	389A	14490
x"00",	-- Hex Addr	389B	14491
x"00",	-- Hex Addr	389C	14492
x"00",	-- Hex Addr	389D	14493
x"00",	-- Hex Addr	389E	14494
x"00",	-- Hex Addr	389F	14495
x"00",	-- Hex Addr	38A0	14496
x"00",	-- Hex Addr	38A1	14497
x"00",	-- Hex Addr	38A2	14498
x"00",	-- Hex Addr	38A3	14499
x"00",	-- Hex Addr	38A4	14500
x"00",	-- Hex Addr	38A5	14501
x"00",	-- Hex Addr	38A6	14502
x"00",	-- Hex Addr	38A7	14503
x"00",	-- Hex Addr	38A8	14504
x"00",	-- Hex Addr	38A9	14505
x"00",	-- Hex Addr	38AA	14506
x"00",	-- Hex Addr	38AB	14507
x"00",	-- Hex Addr	38AC	14508
x"00",	-- Hex Addr	38AD	14509
x"00",	-- Hex Addr	38AE	14510
x"00",	-- Hex Addr	38AF	14511
x"00",	-- Hex Addr	38B0	14512
x"00",	-- Hex Addr	38B1	14513
x"00",	-- Hex Addr	38B2	14514
x"00",	-- Hex Addr	38B3	14515
x"00",	-- Hex Addr	38B4	14516
x"00",	-- Hex Addr	38B5	14517
x"00",	-- Hex Addr	38B6	14518
x"00",	-- Hex Addr	38B7	14519
x"00",	-- Hex Addr	38B8	14520
x"00",	-- Hex Addr	38B9	14521
x"00",	-- Hex Addr	38BA	14522
x"00",	-- Hex Addr	38BB	14523
x"00",	-- Hex Addr	38BC	14524
x"00",	-- Hex Addr	38BD	14525
x"00",	-- Hex Addr	38BE	14526
x"00",	-- Hex Addr	38BF	14527
x"00",	-- Hex Addr	38C0	14528
x"00",	-- Hex Addr	38C1	14529
x"00",	-- Hex Addr	38C2	14530
x"00",	-- Hex Addr	38C3	14531
x"00",	-- Hex Addr	38C4	14532
x"00",	-- Hex Addr	38C5	14533
x"00",	-- Hex Addr	38C6	14534
x"00",	-- Hex Addr	38C7	14535
x"00",	-- Hex Addr	38C8	14536
x"00",	-- Hex Addr	38C9	14537
x"00",	-- Hex Addr	38CA	14538
x"00",	-- Hex Addr	38CB	14539
x"00",	-- Hex Addr	38CC	14540
x"00",	-- Hex Addr	38CD	14541
x"00",	-- Hex Addr	38CE	14542
x"00",	-- Hex Addr	38CF	14543
x"00",	-- Hex Addr	38D0	14544
x"00",	-- Hex Addr	38D1	14545
x"00",	-- Hex Addr	38D2	14546
x"00",	-- Hex Addr	38D3	14547
x"00",	-- Hex Addr	38D4	14548
x"00",	-- Hex Addr	38D5	14549
x"00",	-- Hex Addr	38D6	14550
x"00",	-- Hex Addr	38D7	14551
x"00",	-- Hex Addr	38D8	14552
x"00",	-- Hex Addr	38D9	14553
x"00",	-- Hex Addr	38DA	14554
x"00",	-- Hex Addr	38DB	14555
x"00",	-- Hex Addr	38DC	14556
x"00",	-- Hex Addr	38DD	14557
x"00",	-- Hex Addr	38DE	14558
x"00",	-- Hex Addr	38DF	14559
x"00",	-- Hex Addr	38E0	14560
x"00",	-- Hex Addr	38E1	14561
x"00",	-- Hex Addr	38E2	14562
x"00",	-- Hex Addr	38E3	14563
x"00",	-- Hex Addr	38E4	14564
x"00",	-- Hex Addr	38E5	14565
x"00",	-- Hex Addr	38E6	14566
x"00",	-- Hex Addr	38E7	14567
x"00",	-- Hex Addr	38E8	14568
x"00",	-- Hex Addr	38E9	14569
x"00",	-- Hex Addr	38EA	14570
x"00",	-- Hex Addr	38EB	14571
x"00",	-- Hex Addr	38EC	14572
x"00",	-- Hex Addr	38ED	14573
x"00",	-- Hex Addr	38EE	14574
x"00",	-- Hex Addr	38EF	14575
x"00",	-- Hex Addr	38F0	14576
x"00",	-- Hex Addr	38F1	14577
x"00",	-- Hex Addr	38F2	14578
x"00",	-- Hex Addr	38F3	14579
x"00",	-- Hex Addr	38F4	14580
x"00",	-- Hex Addr	38F5	14581
x"00",	-- Hex Addr	38F6	14582
x"00",	-- Hex Addr	38F7	14583
x"00",	-- Hex Addr	38F8	14584
x"00",	-- Hex Addr	38F9	14585
x"00",	-- Hex Addr	38FA	14586
x"00",	-- Hex Addr	38FB	14587
x"00",	-- Hex Addr	38FC	14588
x"00",	-- Hex Addr	38FD	14589
x"00",	-- Hex Addr	38FE	14590
x"00",	-- Hex Addr	38FF	14591
x"00",	-- Hex Addr	3900	14592
x"00",	-- Hex Addr	3901	14593
x"00",	-- Hex Addr	3902	14594
x"00",	-- Hex Addr	3903	14595
x"00",	-- Hex Addr	3904	14596
x"00",	-- Hex Addr	3905	14597
x"00",	-- Hex Addr	3906	14598
x"00",	-- Hex Addr	3907	14599
x"00",	-- Hex Addr	3908	14600
x"00",	-- Hex Addr	3909	14601
x"00",	-- Hex Addr	390A	14602
x"00",	-- Hex Addr	390B	14603
x"00",	-- Hex Addr	390C	14604
x"00",	-- Hex Addr	390D	14605
x"00",	-- Hex Addr	390E	14606
x"00",	-- Hex Addr	390F	14607
x"00",	-- Hex Addr	3910	14608
x"00",	-- Hex Addr	3911	14609
x"00",	-- Hex Addr	3912	14610
x"00",	-- Hex Addr	3913	14611
x"00",	-- Hex Addr	3914	14612
x"00",	-- Hex Addr	3915	14613
x"00",	-- Hex Addr	3916	14614
x"00",	-- Hex Addr	3917	14615
x"00",	-- Hex Addr	3918	14616
x"00",	-- Hex Addr	3919	14617
x"00",	-- Hex Addr	391A	14618
x"00",	-- Hex Addr	391B	14619
x"00",	-- Hex Addr	391C	14620
x"00",	-- Hex Addr	391D	14621
x"00",	-- Hex Addr	391E	14622
x"00",	-- Hex Addr	391F	14623
x"00",	-- Hex Addr	3920	14624
x"00",	-- Hex Addr	3921	14625
x"00",	-- Hex Addr	3922	14626
x"00",	-- Hex Addr	3923	14627
x"00",	-- Hex Addr	3924	14628
x"00",	-- Hex Addr	3925	14629
x"00",	-- Hex Addr	3926	14630
x"00",	-- Hex Addr	3927	14631
x"00",	-- Hex Addr	3928	14632
x"00",	-- Hex Addr	3929	14633
x"00",	-- Hex Addr	392A	14634
x"00",	-- Hex Addr	392B	14635
x"00",	-- Hex Addr	392C	14636
x"00",	-- Hex Addr	392D	14637
x"00",	-- Hex Addr	392E	14638
x"00",	-- Hex Addr	392F	14639
x"00",	-- Hex Addr	3930	14640
x"00",	-- Hex Addr	3931	14641
x"00",	-- Hex Addr	3932	14642
x"00",	-- Hex Addr	3933	14643
x"00",	-- Hex Addr	3934	14644
x"00",	-- Hex Addr	3935	14645
x"00",	-- Hex Addr	3936	14646
x"00",	-- Hex Addr	3937	14647
x"00",	-- Hex Addr	3938	14648
x"00",	-- Hex Addr	3939	14649
x"00",	-- Hex Addr	393A	14650
x"00",	-- Hex Addr	393B	14651
x"00",	-- Hex Addr	393C	14652
x"00",	-- Hex Addr	393D	14653
x"00",	-- Hex Addr	393E	14654
x"00",	-- Hex Addr	393F	14655
x"00",	-- Hex Addr	3940	14656
x"00",	-- Hex Addr	3941	14657
x"00",	-- Hex Addr	3942	14658
x"00",	-- Hex Addr	3943	14659
x"00",	-- Hex Addr	3944	14660
x"00",	-- Hex Addr	3945	14661
x"00",	-- Hex Addr	3946	14662
x"00",	-- Hex Addr	3947	14663
x"00",	-- Hex Addr	3948	14664
x"00",	-- Hex Addr	3949	14665
x"00",	-- Hex Addr	394A	14666
x"00",	-- Hex Addr	394B	14667
x"00",	-- Hex Addr	394C	14668
x"00",	-- Hex Addr	394D	14669
x"00",	-- Hex Addr	394E	14670
x"00",	-- Hex Addr	394F	14671
x"00",	-- Hex Addr	3950	14672
x"00",	-- Hex Addr	3951	14673
x"00",	-- Hex Addr	3952	14674
x"00",	-- Hex Addr	3953	14675
x"00",	-- Hex Addr	3954	14676
x"00",	-- Hex Addr	3955	14677
x"00",	-- Hex Addr	3956	14678
x"00",	-- Hex Addr	3957	14679
x"00",	-- Hex Addr	3958	14680
x"00",	-- Hex Addr	3959	14681
x"00",	-- Hex Addr	395A	14682
x"00",	-- Hex Addr	395B	14683
x"00",	-- Hex Addr	395C	14684
x"00",	-- Hex Addr	395D	14685
x"00",	-- Hex Addr	395E	14686
x"00",	-- Hex Addr	395F	14687
x"00",	-- Hex Addr	3960	14688
x"00",	-- Hex Addr	3961	14689
x"00",	-- Hex Addr	3962	14690
x"00",	-- Hex Addr	3963	14691
x"00",	-- Hex Addr	3964	14692
x"00",	-- Hex Addr	3965	14693
x"00",	-- Hex Addr	3966	14694
x"00",	-- Hex Addr	3967	14695
x"00",	-- Hex Addr	3968	14696
x"00",	-- Hex Addr	3969	14697
x"00",	-- Hex Addr	396A	14698
x"00",	-- Hex Addr	396B	14699
x"00",	-- Hex Addr	396C	14700
x"00",	-- Hex Addr	396D	14701
x"00",	-- Hex Addr	396E	14702
x"00",	-- Hex Addr	396F	14703
x"00",	-- Hex Addr	3970	14704
x"00",	-- Hex Addr	3971	14705
x"00",	-- Hex Addr	3972	14706
x"00",	-- Hex Addr	3973	14707
x"00",	-- Hex Addr	3974	14708
x"00",	-- Hex Addr	3975	14709
x"00",	-- Hex Addr	3976	14710
x"00",	-- Hex Addr	3977	14711
x"00",	-- Hex Addr	3978	14712
x"00",	-- Hex Addr	3979	14713
x"00",	-- Hex Addr	397A	14714
x"00",	-- Hex Addr	397B	14715
x"00",	-- Hex Addr	397C	14716
x"00",	-- Hex Addr	397D	14717
x"00",	-- Hex Addr	397E	14718
x"00",	-- Hex Addr	397F	14719
x"00",	-- Hex Addr	3980	14720
x"00",	-- Hex Addr	3981	14721
x"00",	-- Hex Addr	3982	14722
x"00",	-- Hex Addr	3983	14723
x"00",	-- Hex Addr	3984	14724
x"00",	-- Hex Addr	3985	14725
x"00",	-- Hex Addr	3986	14726
x"00",	-- Hex Addr	3987	14727
x"00",	-- Hex Addr	3988	14728
x"00",	-- Hex Addr	3989	14729
x"00",	-- Hex Addr	398A	14730
x"00",	-- Hex Addr	398B	14731
x"00",	-- Hex Addr	398C	14732
x"00",	-- Hex Addr	398D	14733
x"00",	-- Hex Addr	398E	14734
x"00",	-- Hex Addr	398F	14735
x"00",	-- Hex Addr	3990	14736
x"00",	-- Hex Addr	3991	14737
x"00",	-- Hex Addr	3992	14738
x"00",	-- Hex Addr	3993	14739
x"00",	-- Hex Addr	3994	14740
x"00",	-- Hex Addr	3995	14741
x"00",	-- Hex Addr	3996	14742
x"00",	-- Hex Addr	3997	14743
x"00",	-- Hex Addr	3998	14744
x"00",	-- Hex Addr	3999	14745
x"00",	-- Hex Addr	399A	14746
x"00",	-- Hex Addr	399B	14747
x"00",	-- Hex Addr	399C	14748
x"00",	-- Hex Addr	399D	14749
x"00",	-- Hex Addr	399E	14750
x"00",	-- Hex Addr	399F	14751
x"00",	-- Hex Addr	39A0	14752
x"00",	-- Hex Addr	39A1	14753
x"00",	-- Hex Addr	39A2	14754
x"00",	-- Hex Addr	39A3	14755
x"00",	-- Hex Addr	39A4	14756
x"00",	-- Hex Addr	39A5	14757
x"00",	-- Hex Addr	39A6	14758
x"00",	-- Hex Addr	39A7	14759
x"00",	-- Hex Addr	39A8	14760
x"00",	-- Hex Addr	39A9	14761
x"00",	-- Hex Addr	39AA	14762
x"00",	-- Hex Addr	39AB	14763
x"00",	-- Hex Addr	39AC	14764
x"00",	-- Hex Addr	39AD	14765
x"00",	-- Hex Addr	39AE	14766
x"00",	-- Hex Addr	39AF	14767
x"00",	-- Hex Addr	39B0	14768
x"00",	-- Hex Addr	39B1	14769
x"00",	-- Hex Addr	39B2	14770
x"00",	-- Hex Addr	39B3	14771
x"00",	-- Hex Addr	39B4	14772
x"00",	-- Hex Addr	39B5	14773
x"00",	-- Hex Addr	39B6	14774
x"00",	-- Hex Addr	39B7	14775
x"00",	-- Hex Addr	39B8	14776
x"00",	-- Hex Addr	39B9	14777
x"00",	-- Hex Addr	39BA	14778
x"00",	-- Hex Addr	39BB	14779
x"00",	-- Hex Addr	39BC	14780
x"00",	-- Hex Addr	39BD	14781
x"00",	-- Hex Addr	39BE	14782
x"00",	-- Hex Addr	39BF	14783
x"00",	-- Hex Addr	39C0	14784
x"00",	-- Hex Addr	39C1	14785
x"00",	-- Hex Addr	39C2	14786
x"00",	-- Hex Addr	39C3	14787
x"00",	-- Hex Addr	39C4	14788
x"00",	-- Hex Addr	39C5	14789
x"00",	-- Hex Addr	39C6	14790
x"00",	-- Hex Addr	39C7	14791
x"00",	-- Hex Addr	39C8	14792
x"00",	-- Hex Addr	39C9	14793
x"00",	-- Hex Addr	39CA	14794
x"00",	-- Hex Addr	39CB	14795
x"00",	-- Hex Addr	39CC	14796
x"00",	-- Hex Addr	39CD	14797
x"00",	-- Hex Addr	39CE	14798
x"00",	-- Hex Addr	39CF	14799
x"00",	-- Hex Addr	39D0	14800
x"00",	-- Hex Addr	39D1	14801
x"00",	-- Hex Addr	39D2	14802
x"00",	-- Hex Addr	39D3	14803
x"00",	-- Hex Addr	39D4	14804
x"00",	-- Hex Addr	39D5	14805
x"00",	-- Hex Addr	39D6	14806
x"00",	-- Hex Addr	39D7	14807
x"00",	-- Hex Addr	39D8	14808
x"00",	-- Hex Addr	39D9	14809
x"00",	-- Hex Addr	39DA	14810
x"00",	-- Hex Addr	39DB	14811
x"00",	-- Hex Addr	39DC	14812
x"00",	-- Hex Addr	39DD	14813
x"00",	-- Hex Addr	39DE	14814
x"00",	-- Hex Addr	39DF	14815
x"00",	-- Hex Addr	39E0	14816
x"00",	-- Hex Addr	39E1	14817
x"00",	-- Hex Addr	39E2	14818
x"00",	-- Hex Addr	39E3	14819
x"00",	-- Hex Addr	39E4	14820
x"00",	-- Hex Addr	39E5	14821
x"00",	-- Hex Addr	39E6	14822
x"00",	-- Hex Addr	39E7	14823
x"00",	-- Hex Addr	39E8	14824
x"00",	-- Hex Addr	39E9	14825
x"00",	-- Hex Addr	39EA	14826
x"00",	-- Hex Addr	39EB	14827
x"00",	-- Hex Addr	39EC	14828
x"00",	-- Hex Addr	39ED	14829
x"00",	-- Hex Addr	39EE	14830
x"00",	-- Hex Addr	39EF	14831
x"00",	-- Hex Addr	39F0	14832
x"00",	-- Hex Addr	39F1	14833
x"00",	-- Hex Addr	39F2	14834
x"00",	-- Hex Addr	39F3	14835
x"00",	-- Hex Addr	39F4	14836
x"00",	-- Hex Addr	39F5	14837
x"00",	-- Hex Addr	39F6	14838
x"00",	-- Hex Addr	39F7	14839
x"00",	-- Hex Addr	39F8	14840
x"00",	-- Hex Addr	39F9	14841
x"00",	-- Hex Addr	39FA	14842
x"00",	-- Hex Addr	39FB	14843
x"00",	-- Hex Addr	39FC	14844
x"00",	-- Hex Addr	39FD	14845
x"00",	-- Hex Addr	39FE	14846
x"00",	-- Hex Addr	39FF	14847
x"00",	-- Hex Addr	3A00	14848
x"00",	-- Hex Addr	3A01	14849
x"00",	-- Hex Addr	3A02	14850
x"00",	-- Hex Addr	3A03	14851
x"00",	-- Hex Addr	3A04	14852
x"00",	-- Hex Addr	3A05	14853
x"00",	-- Hex Addr	3A06	14854
x"00",	-- Hex Addr	3A07	14855
x"00",	-- Hex Addr	3A08	14856
x"00",	-- Hex Addr	3A09	14857
x"00",	-- Hex Addr	3A0A	14858
x"00",	-- Hex Addr	3A0B	14859
x"00",	-- Hex Addr	3A0C	14860
x"00",	-- Hex Addr	3A0D	14861
x"00",	-- Hex Addr	3A0E	14862
x"00",	-- Hex Addr	3A0F	14863
x"00",	-- Hex Addr	3A10	14864
x"00",	-- Hex Addr	3A11	14865
x"00",	-- Hex Addr	3A12	14866
x"00",	-- Hex Addr	3A13	14867
x"00",	-- Hex Addr	3A14	14868
x"00",	-- Hex Addr	3A15	14869
x"00",	-- Hex Addr	3A16	14870
x"00",	-- Hex Addr	3A17	14871
x"00",	-- Hex Addr	3A18	14872
x"00",	-- Hex Addr	3A19	14873
x"00",	-- Hex Addr	3A1A	14874
x"00",	-- Hex Addr	3A1B	14875
x"00",	-- Hex Addr	3A1C	14876
x"00",	-- Hex Addr	3A1D	14877
x"00",	-- Hex Addr	3A1E	14878
x"00",	-- Hex Addr	3A1F	14879
x"00",	-- Hex Addr	3A20	14880
x"00",	-- Hex Addr	3A21	14881
x"00",	-- Hex Addr	3A22	14882
x"00",	-- Hex Addr	3A23	14883
x"00",	-- Hex Addr	3A24	14884
x"00",	-- Hex Addr	3A25	14885
x"00",	-- Hex Addr	3A26	14886
x"00",	-- Hex Addr	3A27	14887
x"00",	-- Hex Addr	3A28	14888
x"00",	-- Hex Addr	3A29	14889
x"00",	-- Hex Addr	3A2A	14890
x"00",	-- Hex Addr	3A2B	14891
x"00",	-- Hex Addr	3A2C	14892
x"00",	-- Hex Addr	3A2D	14893
x"00",	-- Hex Addr	3A2E	14894
x"00",	-- Hex Addr	3A2F	14895
x"00",	-- Hex Addr	3A30	14896
x"00",	-- Hex Addr	3A31	14897
x"00",	-- Hex Addr	3A32	14898
x"00",	-- Hex Addr	3A33	14899
x"00",	-- Hex Addr	3A34	14900
x"00",	-- Hex Addr	3A35	14901
x"00",	-- Hex Addr	3A36	14902
x"00",	-- Hex Addr	3A37	14903
x"00",	-- Hex Addr	3A38	14904
x"00",	-- Hex Addr	3A39	14905
x"00",	-- Hex Addr	3A3A	14906
x"00",	-- Hex Addr	3A3B	14907
x"00",	-- Hex Addr	3A3C	14908
x"00",	-- Hex Addr	3A3D	14909
x"00",	-- Hex Addr	3A3E	14910
x"00",	-- Hex Addr	3A3F	14911
x"00",	-- Hex Addr	3A40	14912
x"00",	-- Hex Addr	3A41	14913
x"00",	-- Hex Addr	3A42	14914
x"00",	-- Hex Addr	3A43	14915
x"00",	-- Hex Addr	3A44	14916
x"00",	-- Hex Addr	3A45	14917
x"00",	-- Hex Addr	3A46	14918
x"00",	-- Hex Addr	3A47	14919
x"00",	-- Hex Addr	3A48	14920
x"00",	-- Hex Addr	3A49	14921
x"00",	-- Hex Addr	3A4A	14922
x"00",	-- Hex Addr	3A4B	14923
x"00",	-- Hex Addr	3A4C	14924
x"00",	-- Hex Addr	3A4D	14925
x"00",	-- Hex Addr	3A4E	14926
x"00",	-- Hex Addr	3A4F	14927
x"00",	-- Hex Addr	3A50	14928
x"00",	-- Hex Addr	3A51	14929
x"00",	-- Hex Addr	3A52	14930
x"00",	-- Hex Addr	3A53	14931
x"00",	-- Hex Addr	3A54	14932
x"00",	-- Hex Addr	3A55	14933
x"00",	-- Hex Addr	3A56	14934
x"00",	-- Hex Addr	3A57	14935
x"00",	-- Hex Addr	3A58	14936
x"00",	-- Hex Addr	3A59	14937
x"00",	-- Hex Addr	3A5A	14938
x"00",	-- Hex Addr	3A5B	14939
x"00",	-- Hex Addr	3A5C	14940
x"00",	-- Hex Addr	3A5D	14941
x"00",	-- Hex Addr	3A5E	14942
x"00",	-- Hex Addr	3A5F	14943
x"00",	-- Hex Addr	3A60	14944
x"00",	-- Hex Addr	3A61	14945
x"00",	-- Hex Addr	3A62	14946
x"00",	-- Hex Addr	3A63	14947
x"00",	-- Hex Addr	3A64	14948
x"00",	-- Hex Addr	3A65	14949
x"00",	-- Hex Addr	3A66	14950
x"00",	-- Hex Addr	3A67	14951
x"00",	-- Hex Addr	3A68	14952
x"00",	-- Hex Addr	3A69	14953
x"00",	-- Hex Addr	3A6A	14954
x"00",	-- Hex Addr	3A6B	14955
x"00",	-- Hex Addr	3A6C	14956
x"00",	-- Hex Addr	3A6D	14957
x"00",	-- Hex Addr	3A6E	14958
x"00",	-- Hex Addr	3A6F	14959
x"00",	-- Hex Addr	3A70	14960
x"00",	-- Hex Addr	3A71	14961
x"00",	-- Hex Addr	3A72	14962
x"00",	-- Hex Addr	3A73	14963
x"00",	-- Hex Addr	3A74	14964
x"00",	-- Hex Addr	3A75	14965
x"00",	-- Hex Addr	3A76	14966
x"00",	-- Hex Addr	3A77	14967
x"00",	-- Hex Addr	3A78	14968
x"00",	-- Hex Addr	3A79	14969
x"00",	-- Hex Addr	3A7A	14970
x"00",	-- Hex Addr	3A7B	14971
x"00",	-- Hex Addr	3A7C	14972
x"00",	-- Hex Addr	3A7D	14973
x"00",	-- Hex Addr	3A7E	14974
x"00",	-- Hex Addr	3A7F	14975
x"00",	-- Hex Addr	3A80	14976
x"00",	-- Hex Addr	3A81	14977
x"00",	-- Hex Addr	3A82	14978
x"00",	-- Hex Addr	3A83	14979
x"00",	-- Hex Addr	3A84	14980
x"00",	-- Hex Addr	3A85	14981
x"00",	-- Hex Addr	3A86	14982
x"00",	-- Hex Addr	3A87	14983
x"00",	-- Hex Addr	3A88	14984
x"00",	-- Hex Addr	3A89	14985
x"00",	-- Hex Addr	3A8A	14986
x"00",	-- Hex Addr	3A8B	14987
x"00",	-- Hex Addr	3A8C	14988
x"00",	-- Hex Addr	3A8D	14989
x"00",	-- Hex Addr	3A8E	14990
x"00",	-- Hex Addr	3A8F	14991
x"00",	-- Hex Addr	3A90	14992
x"00",	-- Hex Addr	3A91	14993
x"00",	-- Hex Addr	3A92	14994
x"00",	-- Hex Addr	3A93	14995
x"00",	-- Hex Addr	3A94	14996
x"00",	-- Hex Addr	3A95	14997
x"00",	-- Hex Addr	3A96	14998
x"00",	-- Hex Addr	3A97	14999
x"00",	-- Hex Addr	3A98	15000
x"00",	-- Hex Addr	3A99	15001
x"00",	-- Hex Addr	3A9A	15002
x"00",	-- Hex Addr	3A9B	15003
x"00",	-- Hex Addr	3A9C	15004
x"00",	-- Hex Addr	3A9D	15005
x"00",	-- Hex Addr	3A9E	15006
x"00",	-- Hex Addr	3A9F	15007
x"00",	-- Hex Addr	3AA0	15008
x"00",	-- Hex Addr	3AA1	15009
x"00",	-- Hex Addr	3AA2	15010
x"00",	-- Hex Addr	3AA3	15011
x"00",	-- Hex Addr	3AA4	15012
x"00",	-- Hex Addr	3AA5	15013
x"00",	-- Hex Addr	3AA6	15014
x"00",	-- Hex Addr	3AA7	15015
x"00",	-- Hex Addr	3AA8	15016
x"00",	-- Hex Addr	3AA9	15017
x"00",	-- Hex Addr	3AAA	15018
x"00",	-- Hex Addr	3AAB	15019
x"00",	-- Hex Addr	3AAC	15020
x"00",	-- Hex Addr	3AAD	15021
x"00",	-- Hex Addr	3AAE	15022
x"00",	-- Hex Addr	3AAF	15023
x"00",	-- Hex Addr	3AB0	15024
x"00",	-- Hex Addr	3AB1	15025
x"00",	-- Hex Addr	3AB2	15026
x"00",	-- Hex Addr	3AB3	15027
x"00",	-- Hex Addr	3AB4	15028
x"00",	-- Hex Addr	3AB5	15029
x"00",	-- Hex Addr	3AB6	15030
x"00",	-- Hex Addr	3AB7	15031
x"00",	-- Hex Addr	3AB8	15032
x"00",	-- Hex Addr	3AB9	15033
x"00",	-- Hex Addr	3ABA	15034
x"00",	-- Hex Addr	3ABB	15035
x"00",	-- Hex Addr	3ABC	15036
x"00",	-- Hex Addr	3ABD	15037
x"00",	-- Hex Addr	3ABE	15038
x"00",	-- Hex Addr	3ABF	15039
x"00",	-- Hex Addr	3AC0	15040
x"00",	-- Hex Addr	3AC1	15041
x"00",	-- Hex Addr	3AC2	15042
x"00",	-- Hex Addr	3AC3	15043
x"00",	-- Hex Addr	3AC4	15044
x"00",	-- Hex Addr	3AC5	15045
x"00",	-- Hex Addr	3AC6	15046
x"00",	-- Hex Addr	3AC7	15047
x"00",	-- Hex Addr	3AC8	15048
x"00",	-- Hex Addr	3AC9	15049
x"00",	-- Hex Addr	3ACA	15050
x"00",	-- Hex Addr	3ACB	15051
x"00",	-- Hex Addr	3ACC	15052
x"00",	-- Hex Addr	3ACD	15053
x"00",	-- Hex Addr	3ACE	15054
x"00",	-- Hex Addr	3ACF	15055
x"00",	-- Hex Addr	3AD0	15056
x"00",	-- Hex Addr	3AD1	15057
x"00",	-- Hex Addr	3AD2	15058
x"00",	-- Hex Addr	3AD3	15059
x"00",	-- Hex Addr	3AD4	15060
x"00",	-- Hex Addr	3AD5	15061
x"00",	-- Hex Addr	3AD6	15062
x"00",	-- Hex Addr	3AD7	15063
x"00",	-- Hex Addr	3AD8	15064
x"00",	-- Hex Addr	3AD9	15065
x"00",	-- Hex Addr	3ADA	15066
x"00",	-- Hex Addr	3ADB	15067
x"00",	-- Hex Addr	3ADC	15068
x"00",	-- Hex Addr	3ADD	15069
x"00",	-- Hex Addr	3ADE	15070
x"00",	-- Hex Addr	3ADF	15071
x"00",	-- Hex Addr	3AE0	15072
x"00",	-- Hex Addr	3AE1	15073
x"00",	-- Hex Addr	3AE2	15074
x"00",	-- Hex Addr	3AE3	15075
x"00",	-- Hex Addr	3AE4	15076
x"00",	-- Hex Addr	3AE5	15077
x"00",	-- Hex Addr	3AE6	15078
x"00",	-- Hex Addr	3AE7	15079
x"00",	-- Hex Addr	3AE8	15080
x"00",	-- Hex Addr	3AE9	15081
x"00",	-- Hex Addr	3AEA	15082
x"00",	-- Hex Addr	3AEB	15083
x"00",	-- Hex Addr	3AEC	15084
x"00",	-- Hex Addr	3AED	15085
x"00",	-- Hex Addr	3AEE	15086
x"00",	-- Hex Addr	3AEF	15087
x"00",	-- Hex Addr	3AF0	15088
x"00",	-- Hex Addr	3AF1	15089
x"00",	-- Hex Addr	3AF2	15090
x"00",	-- Hex Addr	3AF3	15091
x"00",	-- Hex Addr	3AF4	15092
x"00",	-- Hex Addr	3AF5	15093
x"00",	-- Hex Addr	3AF6	15094
x"00",	-- Hex Addr	3AF7	15095
x"00",	-- Hex Addr	3AF8	15096
x"00",	-- Hex Addr	3AF9	15097
x"00",	-- Hex Addr	3AFA	15098
x"00",	-- Hex Addr	3AFB	15099
x"00",	-- Hex Addr	3AFC	15100
x"00",	-- Hex Addr	3AFD	15101
x"00",	-- Hex Addr	3AFE	15102
x"00",	-- Hex Addr	3AFF	15103
x"00",	-- Hex Addr	3B00	15104
x"00",	-- Hex Addr	3B01	15105
x"00",	-- Hex Addr	3B02	15106
x"00",	-- Hex Addr	3B03	15107
x"00",	-- Hex Addr	3B04	15108
x"00",	-- Hex Addr	3B05	15109
x"00",	-- Hex Addr	3B06	15110
x"00",	-- Hex Addr	3B07	15111
x"00",	-- Hex Addr	3B08	15112
x"00",	-- Hex Addr	3B09	15113
x"00",	-- Hex Addr	3B0A	15114
x"00",	-- Hex Addr	3B0B	15115
x"00",	-- Hex Addr	3B0C	15116
x"00",	-- Hex Addr	3B0D	15117
x"00",	-- Hex Addr	3B0E	15118
x"00",	-- Hex Addr	3B0F	15119
x"00",	-- Hex Addr	3B10	15120
x"00",	-- Hex Addr	3B11	15121
x"00",	-- Hex Addr	3B12	15122
x"00",	-- Hex Addr	3B13	15123
x"00",	-- Hex Addr	3B14	15124
x"00",	-- Hex Addr	3B15	15125
x"00",	-- Hex Addr	3B16	15126
x"00",	-- Hex Addr	3B17	15127
x"00",	-- Hex Addr	3B18	15128
x"00",	-- Hex Addr	3B19	15129
x"00",	-- Hex Addr	3B1A	15130
x"00",	-- Hex Addr	3B1B	15131
x"00",	-- Hex Addr	3B1C	15132
x"00",	-- Hex Addr	3B1D	15133
x"00",	-- Hex Addr	3B1E	15134
x"00",	-- Hex Addr	3B1F	15135
x"00",	-- Hex Addr	3B20	15136
x"00",	-- Hex Addr	3B21	15137
x"00",	-- Hex Addr	3B22	15138
x"00",	-- Hex Addr	3B23	15139
x"00",	-- Hex Addr	3B24	15140
x"00",	-- Hex Addr	3B25	15141
x"00",	-- Hex Addr	3B26	15142
x"00",	-- Hex Addr	3B27	15143
x"00",	-- Hex Addr	3B28	15144
x"00",	-- Hex Addr	3B29	15145
x"00",	-- Hex Addr	3B2A	15146
x"00",	-- Hex Addr	3B2B	15147
x"00",	-- Hex Addr	3B2C	15148
x"00",	-- Hex Addr	3B2D	15149
x"00",	-- Hex Addr	3B2E	15150
x"00",	-- Hex Addr	3B2F	15151
x"00",	-- Hex Addr	3B30	15152
x"00",	-- Hex Addr	3B31	15153
x"00",	-- Hex Addr	3B32	15154
x"00",	-- Hex Addr	3B33	15155
x"00",	-- Hex Addr	3B34	15156
x"00",	-- Hex Addr	3B35	15157
x"00",	-- Hex Addr	3B36	15158
x"00",	-- Hex Addr	3B37	15159
x"00",	-- Hex Addr	3B38	15160
x"00",	-- Hex Addr	3B39	15161
x"00",	-- Hex Addr	3B3A	15162
x"00",	-- Hex Addr	3B3B	15163
x"00",	-- Hex Addr	3B3C	15164
x"00",	-- Hex Addr	3B3D	15165
x"00",	-- Hex Addr	3B3E	15166
x"00",	-- Hex Addr	3B3F	15167
x"00",	-- Hex Addr	3B40	15168
x"00",	-- Hex Addr	3B41	15169
x"00",	-- Hex Addr	3B42	15170
x"00",	-- Hex Addr	3B43	15171
x"00",	-- Hex Addr	3B44	15172
x"00",	-- Hex Addr	3B45	15173
x"00",	-- Hex Addr	3B46	15174
x"00",	-- Hex Addr	3B47	15175
x"00",	-- Hex Addr	3B48	15176
x"00",	-- Hex Addr	3B49	15177
x"00",	-- Hex Addr	3B4A	15178
x"00",	-- Hex Addr	3B4B	15179
x"00",	-- Hex Addr	3B4C	15180
x"00",	-- Hex Addr	3B4D	15181
x"00",	-- Hex Addr	3B4E	15182
x"00",	-- Hex Addr	3B4F	15183
x"00",	-- Hex Addr	3B50	15184
x"00",	-- Hex Addr	3B51	15185
x"00",	-- Hex Addr	3B52	15186
x"00",	-- Hex Addr	3B53	15187
x"00",	-- Hex Addr	3B54	15188
x"00",	-- Hex Addr	3B55	15189
x"00",	-- Hex Addr	3B56	15190
x"00",	-- Hex Addr	3B57	15191
x"00",	-- Hex Addr	3B58	15192
x"00",	-- Hex Addr	3B59	15193
x"00",	-- Hex Addr	3B5A	15194
x"00",	-- Hex Addr	3B5B	15195
x"00",	-- Hex Addr	3B5C	15196
x"00",	-- Hex Addr	3B5D	15197
x"00",	-- Hex Addr	3B5E	15198
x"00",	-- Hex Addr	3B5F	15199
x"00",	-- Hex Addr	3B60	15200
x"00",	-- Hex Addr	3B61	15201
x"00",	-- Hex Addr	3B62	15202
x"00",	-- Hex Addr	3B63	15203
x"00",	-- Hex Addr	3B64	15204
x"00",	-- Hex Addr	3B65	15205
x"00",	-- Hex Addr	3B66	15206
x"00",	-- Hex Addr	3B67	15207
x"00",	-- Hex Addr	3B68	15208
x"00",	-- Hex Addr	3B69	15209
x"00",	-- Hex Addr	3B6A	15210
x"00",	-- Hex Addr	3B6B	15211
x"00",	-- Hex Addr	3B6C	15212
x"00",	-- Hex Addr	3B6D	15213
x"00",	-- Hex Addr	3B6E	15214
x"00",	-- Hex Addr	3B6F	15215
x"00",	-- Hex Addr	3B70	15216
x"00",	-- Hex Addr	3B71	15217
x"00",	-- Hex Addr	3B72	15218
x"00",	-- Hex Addr	3B73	15219
x"00",	-- Hex Addr	3B74	15220
x"00",	-- Hex Addr	3B75	15221
x"00",	-- Hex Addr	3B76	15222
x"00",	-- Hex Addr	3B77	15223
x"00",	-- Hex Addr	3B78	15224
x"00",	-- Hex Addr	3B79	15225
x"00",	-- Hex Addr	3B7A	15226
x"00",	-- Hex Addr	3B7B	15227
x"00",	-- Hex Addr	3B7C	15228
x"00",	-- Hex Addr	3B7D	15229
x"00",	-- Hex Addr	3B7E	15230
x"00",	-- Hex Addr	3B7F	15231
x"00",	-- Hex Addr	3B80	15232
x"00",	-- Hex Addr	3B81	15233
x"00",	-- Hex Addr	3B82	15234
x"00",	-- Hex Addr	3B83	15235
x"00",	-- Hex Addr	3B84	15236
x"00",	-- Hex Addr	3B85	15237
x"00",	-- Hex Addr	3B86	15238
x"00",	-- Hex Addr	3B87	15239
x"00",	-- Hex Addr	3B88	15240
x"00",	-- Hex Addr	3B89	15241
x"00",	-- Hex Addr	3B8A	15242
x"00",	-- Hex Addr	3B8B	15243
x"00",	-- Hex Addr	3B8C	15244
x"00",	-- Hex Addr	3B8D	15245
x"00",	-- Hex Addr	3B8E	15246
x"00",	-- Hex Addr	3B8F	15247
x"00",	-- Hex Addr	3B90	15248
x"00",	-- Hex Addr	3B91	15249
x"00",	-- Hex Addr	3B92	15250
x"00",	-- Hex Addr	3B93	15251
x"00",	-- Hex Addr	3B94	15252
x"00",	-- Hex Addr	3B95	15253
x"00",	-- Hex Addr	3B96	15254
x"00",	-- Hex Addr	3B97	15255
x"00",	-- Hex Addr	3B98	15256
x"00",	-- Hex Addr	3B99	15257
x"00",	-- Hex Addr	3B9A	15258
x"00",	-- Hex Addr	3B9B	15259
x"00",	-- Hex Addr	3B9C	15260
x"00",	-- Hex Addr	3B9D	15261
x"00",	-- Hex Addr	3B9E	15262
x"00",	-- Hex Addr	3B9F	15263
x"00",	-- Hex Addr	3BA0	15264
x"00",	-- Hex Addr	3BA1	15265
x"00",	-- Hex Addr	3BA2	15266
x"00",	-- Hex Addr	3BA3	15267
x"00",	-- Hex Addr	3BA4	15268
x"00",	-- Hex Addr	3BA5	15269
x"00",	-- Hex Addr	3BA6	15270
x"00",	-- Hex Addr	3BA7	15271
x"00",	-- Hex Addr	3BA8	15272
x"00",	-- Hex Addr	3BA9	15273
x"00",	-- Hex Addr	3BAA	15274
x"00",	-- Hex Addr	3BAB	15275
x"00",	-- Hex Addr	3BAC	15276
x"00",	-- Hex Addr	3BAD	15277
x"00",	-- Hex Addr	3BAE	15278
x"00",	-- Hex Addr	3BAF	15279
x"00",	-- Hex Addr	3BB0	15280
x"00",	-- Hex Addr	3BB1	15281
x"00",	-- Hex Addr	3BB2	15282
x"00",	-- Hex Addr	3BB3	15283
x"00",	-- Hex Addr	3BB4	15284
x"00",	-- Hex Addr	3BB5	15285
x"00",	-- Hex Addr	3BB6	15286
x"00",	-- Hex Addr	3BB7	15287
x"00",	-- Hex Addr	3BB8	15288
x"00",	-- Hex Addr	3BB9	15289
x"00",	-- Hex Addr	3BBA	15290
x"00",	-- Hex Addr	3BBB	15291
x"00",	-- Hex Addr	3BBC	15292
x"00",	-- Hex Addr	3BBD	15293
x"00",	-- Hex Addr	3BBE	15294
x"00",	-- Hex Addr	3BBF	15295
x"00",	-- Hex Addr	3BC0	15296
x"00",	-- Hex Addr	3BC1	15297
x"00",	-- Hex Addr	3BC2	15298
x"00",	-- Hex Addr	3BC3	15299
x"00",	-- Hex Addr	3BC4	15300
x"00",	-- Hex Addr	3BC5	15301
x"00",	-- Hex Addr	3BC6	15302
x"00",	-- Hex Addr	3BC7	15303
x"00",	-- Hex Addr	3BC8	15304
x"00",	-- Hex Addr	3BC9	15305
x"00",	-- Hex Addr	3BCA	15306
x"00",	-- Hex Addr	3BCB	15307
x"00",	-- Hex Addr	3BCC	15308
x"00",	-- Hex Addr	3BCD	15309
x"00",	-- Hex Addr	3BCE	15310
x"00",	-- Hex Addr	3BCF	15311
x"00",	-- Hex Addr	3BD0	15312
x"00",	-- Hex Addr	3BD1	15313
x"00",	-- Hex Addr	3BD2	15314
x"00",	-- Hex Addr	3BD3	15315
x"00",	-- Hex Addr	3BD4	15316
x"00",	-- Hex Addr	3BD5	15317
x"00",	-- Hex Addr	3BD6	15318
x"00",	-- Hex Addr	3BD7	15319
x"00",	-- Hex Addr	3BD8	15320
x"00",	-- Hex Addr	3BD9	15321
x"00",	-- Hex Addr	3BDA	15322
x"00",	-- Hex Addr	3BDB	15323
x"00",	-- Hex Addr	3BDC	15324
x"00",	-- Hex Addr	3BDD	15325
x"00",	-- Hex Addr	3BDE	15326
x"00",	-- Hex Addr	3BDF	15327
x"00",	-- Hex Addr	3BE0	15328
x"00",	-- Hex Addr	3BE1	15329
x"00",	-- Hex Addr	3BE2	15330
x"00",	-- Hex Addr	3BE3	15331
x"00",	-- Hex Addr	3BE4	15332
x"00",	-- Hex Addr	3BE5	15333
x"00",	-- Hex Addr	3BE6	15334
x"00",	-- Hex Addr	3BE7	15335
x"00",	-- Hex Addr	3BE8	15336
x"00",	-- Hex Addr	3BE9	15337
x"00",	-- Hex Addr	3BEA	15338
x"00",	-- Hex Addr	3BEB	15339
x"00",	-- Hex Addr	3BEC	15340
x"00",	-- Hex Addr	3BED	15341
x"00",	-- Hex Addr	3BEE	15342
x"00",	-- Hex Addr	3BEF	15343
x"00",	-- Hex Addr	3BF0	15344
x"00",	-- Hex Addr	3BF1	15345
x"00",	-- Hex Addr	3BF2	15346
x"00",	-- Hex Addr	3BF3	15347
x"00",	-- Hex Addr	3BF4	15348
x"00",	-- Hex Addr	3BF5	15349
x"00",	-- Hex Addr	3BF6	15350
x"00",	-- Hex Addr	3BF7	15351
x"00",	-- Hex Addr	3BF8	15352
x"00",	-- Hex Addr	3BF9	15353
x"00",	-- Hex Addr	3BFA	15354
x"00",	-- Hex Addr	3BFB	15355
x"00",	-- Hex Addr	3BFC	15356
x"00",	-- Hex Addr	3BFD	15357
x"00",	-- Hex Addr	3BFE	15358
x"00",	-- Hex Addr	3BFF	15359
x"00",	-- Hex Addr	3C00	15360
x"00",	-- Hex Addr	3C01	15361
x"00",	-- Hex Addr	3C02	15362
x"00",	-- Hex Addr	3C03	15363
x"00",	-- Hex Addr	3C04	15364
x"00",	-- Hex Addr	3C05	15365
x"00",	-- Hex Addr	3C06	15366
x"00",	-- Hex Addr	3C07	15367
x"00",	-- Hex Addr	3C08	15368
x"00",	-- Hex Addr	3C09	15369
x"00",	-- Hex Addr	3C0A	15370
x"00",	-- Hex Addr	3C0B	15371
x"00",	-- Hex Addr	3C0C	15372
x"00",	-- Hex Addr	3C0D	15373
x"00",	-- Hex Addr	3C0E	15374
x"00",	-- Hex Addr	3C0F	15375
x"00",	-- Hex Addr	3C10	15376
x"00",	-- Hex Addr	3C11	15377
x"00",	-- Hex Addr	3C12	15378
x"00",	-- Hex Addr	3C13	15379
x"00",	-- Hex Addr	3C14	15380
x"00",	-- Hex Addr	3C15	15381
x"00",	-- Hex Addr	3C16	15382
x"00",	-- Hex Addr	3C17	15383
x"00",	-- Hex Addr	3C18	15384
x"00",	-- Hex Addr	3C19	15385
x"00",	-- Hex Addr	3C1A	15386
x"00",	-- Hex Addr	3C1B	15387
x"00",	-- Hex Addr	3C1C	15388
x"00",	-- Hex Addr	3C1D	15389
x"00",	-- Hex Addr	3C1E	15390
x"00",	-- Hex Addr	3C1F	15391
x"00",	-- Hex Addr	3C20	15392
x"00",	-- Hex Addr	3C21	15393
x"00",	-- Hex Addr	3C22	15394
x"00",	-- Hex Addr	3C23	15395
x"00",	-- Hex Addr	3C24	15396
x"00",	-- Hex Addr	3C25	15397
x"00",	-- Hex Addr	3C26	15398
x"00",	-- Hex Addr	3C27	15399
x"00",	-- Hex Addr	3C28	15400
x"00",	-- Hex Addr	3C29	15401
x"00",	-- Hex Addr	3C2A	15402
x"00",	-- Hex Addr	3C2B	15403
x"00",	-- Hex Addr	3C2C	15404
x"00",	-- Hex Addr	3C2D	15405
x"00",	-- Hex Addr	3C2E	15406
x"00",	-- Hex Addr	3C2F	15407
x"00",	-- Hex Addr	3C30	15408
x"00",	-- Hex Addr	3C31	15409
x"00",	-- Hex Addr	3C32	15410
x"00",	-- Hex Addr	3C33	15411
x"00",	-- Hex Addr	3C34	15412
x"00",	-- Hex Addr	3C35	15413
x"00",	-- Hex Addr	3C36	15414
x"00",	-- Hex Addr	3C37	15415
x"00",	-- Hex Addr	3C38	15416
x"00",	-- Hex Addr	3C39	15417
x"00",	-- Hex Addr	3C3A	15418
x"00",	-- Hex Addr	3C3B	15419
x"00",	-- Hex Addr	3C3C	15420
x"00",	-- Hex Addr	3C3D	15421
x"00",	-- Hex Addr	3C3E	15422
x"00",	-- Hex Addr	3C3F	15423
x"00",	-- Hex Addr	3C40	15424
x"00",	-- Hex Addr	3C41	15425
x"00",	-- Hex Addr	3C42	15426
x"00",	-- Hex Addr	3C43	15427
x"00",	-- Hex Addr	3C44	15428
x"00",	-- Hex Addr	3C45	15429
x"00",	-- Hex Addr	3C46	15430
x"00",	-- Hex Addr	3C47	15431
x"00",	-- Hex Addr	3C48	15432
x"00",	-- Hex Addr	3C49	15433
x"00",	-- Hex Addr	3C4A	15434
x"00",	-- Hex Addr	3C4B	15435
x"00",	-- Hex Addr	3C4C	15436
x"00",	-- Hex Addr	3C4D	15437
x"00",	-- Hex Addr	3C4E	15438
x"00",	-- Hex Addr	3C4F	15439
x"00",	-- Hex Addr	3C50	15440
x"00",	-- Hex Addr	3C51	15441
x"00",	-- Hex Addr	3C52	15442
x"00",	-- Hex Addr	3C53	15443
x"00",	-- Hex Addr	3C54	15444
x"00",	-- Hex Addr	3C55	15445
x"00",	-- Hex Addr	3C56	15446
x"00",	-- Hex Addr	3C57	15447
x"00",	-- Hex Addr	3C58	15448
x"00",	-- Hex Addr	3C59	15449
x"00",	-- Hex Addr	3C5A	15450
x"00",	-- Hex Addr	3C5B	15451
x"00",	-- Hex Addr	3C5C	15452
x"00",	-- Hex Addr	3C5D	15453
x"00",	-- Hex Addr	3C5E	15454
x"00",	-- Hex Addr	3C5F	15455
x"00",	-- Hex Addr	3C60	15456
x"00",	-- Hex Addr	3C61	15457
x"00",	-- Hex Addr	3C62	15458
x"00",	-- Hex Addr	3C63	15459
x"00",	-- Hex Addr	3C64	15460
x"00",	-- Hex Addr	3C65	15461
x"00",	-- Hex Addr	3C66	15462
x"00",	-- Hex Addr	3C67	15463
x"00",	-- Hex Addr	3C68	15464
x"00",	-- Hex Addr	3C69	15465
x"00",	-- Hex Addr	3C6A	15466
x"00",	-- Hex Addr	3C6B	15467
x"00",	-- Hex Addr	3C6C	15468
x"00",	-- Hex Addr	3C6D	15469
x"00",	-- Hex Addr	3C6E	15470
x"00",	-- Hex Addr	3C6F	15471
x"00",	-- Hex Addr	3C70	15472
x"00",	-- Hex Addr	3C71	15473
x"00",	-- Hex Addr	3C72	15474
x"00",	-- Hex Addr	3C73	15475
x"00",	-- Hex Addr	3C74	15476
x"00",	-- Hex Addr	3C75	15477
x"00",	-- Hex Addr	3C76	15478
x"00",	-- Hex Addr	3C77	15479
x"00",	-- Hex Addr	3C78	15480
x"00",	-- Hex Addr	3C79	15481
x"00",	-- Hex Addr	3C7A	15482
x"00",	-- Hex Addr	3C7B	15483
x"00",	-- Hex Addr	3C7C	15484
x"00",	-- Hex Addr	3C7D	15485
x"00",	-- Hex Addr	3C7E	15486
x"00",	-- Hex Addr	3C7F	15487
x"00",	-- Hex Addr	3C80	15488
x"00",	-- Hex Addr	3C81	15489
x"00",	-- Hex Addr	3C82	15490
x"00",	-- Hex Addr	3C83	15491
x"00",	-- Hex Addr	3C84	15492
x"00",	-- Hex Addr	3C85	15493
x"00",	-- Hex Addr	3C86	15494
x"00",	-- Hex Addr	3C87	15495
x"00",	-- Hex Addr	3C88	15496
x"00",	-- Hex Addr	3C89	15497
x"00",	-- Hex Addr	3C8A	15498
x"00",	-- Hex Addr	3C8B	15499
x"00",	-- Hex Addr	3C8C	15500
x"00",	-- Hex Addr	3C8D	15501
x"00",	-- Hex Addr	3C8E	15502
x"00",	-- Hex Addr	3C8F	15503
x"00",	-- Hex Addr	3C90	15504
x"00",	-- Hex Addr	3C91	15505
x"00",	-- Hex Addr	3C92	15506
x"00",	-- Hex Addr	3C93	15507
x"00",	-- Hex Addr	3C94	15508
x"00",	-- Hex Addr	3C95	15509
x"00",	-- Hex Addr	3C96	15510
x"00",	-- Hex Addr	3C97	15511
x"00",	-- Hex Addr	3C98	15512
x"00",	-- Hex Addr	3C99	15513
x"00",	-- Hex Addr	3C9A	15514
x"00",	-- Hex Addr	3C9B	15515
x"00",	-- Hex Addr	3C9C	15516
x"00",	-- Hex Addr	3C9D	15517
x"00",	-- Hex Addr	3C9E	15518
x"00",	-- Hex Addr	3C9F	15519
x"00",	-- Hex Addr	3CA0	15520
x"00",	-- Hex Addr	3CA1	15521
x"00",	-- Hex Addr	3CA2	15522
x"00",	-- Hex Addr	3CA3	15523
x"00",	-- Hex Addr	3CA4	15524
x"00",	-- Hex Addr	3CA5	15525
x"00",	-- Hex Addr	3CA6	15526
x"00",	-- Hex Addr	3CA7	15527
x"00",	-- Hex Addr	3CA8	15528
x"00",	-- Hex Addr	3CA9	15529
x"00",	-- Hex Addr	3CAA	15530
x"00",	-- Hex Addr	3CAB	15531
x"00",	-- Hex Addr	3CAC	15532
x"00",	-- Hex Addr	3CAD	15533
x"00",	-- Hex Addr	3CAE	15534
x"00",	-- Hex Addr	3CAF	15535
x"00",	-- Hex Addr	3CB0	15536
x"00",	-- Hex Addr	3CB1	15537
x"00",	-- Hex Addr	3CB2	15538
x"00",	-- Hex Addr	3CB3	15539
x"00",	-- Hex Addr	3CB4	15540
x"00",	-- Hex Addr	3CB5	15541
x"00",	-- Hex Addr	3CB6	15542
x"00",	-- Hex Addr	3CB7	15543
x"00",	-- Hex Addr	3CB8	15544
x"00",	-- Hex Addr	3CB9	15545
x"00",	-- Hex Addr	3CBA	15546
x"00",	-- Hex Addr	3CBB	15547
x"00",	-- Hex Addr	3CBC	15548
x"00",	-- Hex Addr	3CBD	15549
x"00",	-- Hex Addr	3CBE	15550
x"00",	-- Hex Addr	3CBF	15551
x"00",	-- Hex Addr	3CC0	15552
x"00",	-- Hex Addr	3CC1	15553
x"00",	-- Hex Addr	3CC2	15554
x"00",	-- Hex Addr	3CC3	15555
x"00",	-- Hex Addr	3CC4	15556
x"00",	-- Hex Addr	3CC5	15557
x"00",	-- Hex Addr	3CC6	15558
x"00",	-- Hex Addr	3CC7	15559
x"00",	-- Hex Addr	3CC8	15560
x"00",	-- Hex Addr	3CC9	15561
x"00",	-- Hex Addr	3CCA	15562
x"00",	-- Hex Addr	3CCB	15563
x"00",	-- Hex Addr	3CCC	15564
x"00",	-- Hex Addr	3CCD	15565
x"00",	-- Hex Addr	3CCE	15566
x"00",	-- Hex Addr	3CCF	15567
x"00",	-- Hex Addr	3CD0	15568
x"00",	-- Hex Addr	3CD1	15569
x"00",	-- Hex Addr	3CD2	15570
x"00",	-- Hex Addr	3CD3	15571
x"00",	-- Hex Addr	3CD4	15572
x"00",	-- Hex Addr	3CD5	15573
x"00",	-- Hex Addr	3CD6	15574
x"00",	-- Hex Addr	3CD7	15575
x"00",	-- Hex Addr	3CD8	15576
x"00",	-- Hex Addr	3CD9	15577
x"00",	-- Hex Addr	3CDA	15578
x"00",	-- Hex Addr	3CDB	15579
x"00",	-- Hex Addr	3CDC	15580
x"00",	-- Hex Addr	3CDD	15581
x"00",	-- Hex Addr	3CDE	15582
x"00",	-- Hex Addr	3CDF	15583
x"00",	-- Hex Addr	3CE0	15584
x"00",	-- Hex Addr	3CE1	15585
x"00",	-- Hex Addr	3CE2	15586
x"00",	-- Hex Addr	3CE3	15587
x"00",	-- Hex Addr	3CE4	15588
x"00",	-- Hex Addr	3CE5	15589
x"00",	-- Hex Addr	3CE6	15590
x"00",	-- Hex Addr	3CE7	15591
x"00",	-- Hex Addr	3CE8	15592
x"00",	-- Hex Addr	3CE9	15593
x"00",	-- Hex Addr	3CEA	15594
x"00",	-- Hex Addr	3CEB	15595
x"00",	-- Hex Addr	3CEC	15596
x"00",	-- Hex Addr	3CED	15597
x"00",	-- Hex Addr	3CEE	15598
x"00",	-- Hex Addr	3CEF	15599
x"00",	-- Hex Addr	3CF0	15600
x"00",	-- Hex Addr	3CF1	15601
x"00",	-- Hex Addr	3CF2	15602
x"00",	-- Hex Addr	3CF3	15603
x"00",	-- Hex Addr	3CF4	15604
x"00",	-- Hex Addr	3CF5	15605
x"00",	-- Hex Addr	3CF6	15606
x"00",	-- Hex Addr	3CF7	15607
x"00",	-- Hex Addr	3CF8	15608
x"00",	-- Hex Addr	3CF9	15609
x"00",	-- Hex Addr	3CFA	15610
x"00",	-- Hex Addr	3CFB	15611
x"00",	-- Hex Addr	3CFC	15612
x"00",	-- Hex Addr	3CFD	15613
x"00",	-- Hex Addr	3CFE	15614
x"00",	-- Hex Addr	3CFF	15615
x"00",	-- Hex Addr	3D00	15616
x"00",	-- Hex Addr	3D01	15617
x"00",	-- Hex Addr	3D02	15618
x"00",	-- Hex Addr	3D03	15619
x"00",	-- Hex Addr	3D04	15620
x"00",	-- Hex Addr	3D05	15621
x"00",	-- Hex Addr	3D06	15622
x"00",	-- Hex Addr	3D07	15623
x"00",	-- Hex Addr	3D08	15624
x"00",	-- Hex Addr	3D09	15625
x"00",	-- Hex Addr	3D0A	15626
x"00",	-- Hex Addr	3D0B	15627
x"00",	-- Hex Addr	3D0C	15628
x"00",	-- Hex Addr	3D0D	15629
x"00",	-- Hex Addr	3D0E	15630
x"00",	-- Hex Addr	3D0F	15631
x"00",	-- Hex Addr	3D10	15632
x"00",	-- Hex Addr	3D11	15633
x"00",	-- Hex Addr	3D12	15634
x"00",	-- Hex Addr	3D13	15635
x"00",	-- Hex Addr	3D14	15636
x"00",	-- Hex Addr	3D15	15637
x"00",	-- Hex Addr	3D16	15638
x"00",	-- Hex Addr	3D17	15639
x"00",	-- Hex Addr	3D18	15640
x"00",	-- Hex Addr	3D19	15641
x"00",	-- Hex Addr	3D1A	15642
x"00",	-- Hex Addr	3D1B	15643
x"00",	-- Hex Addr	3D1C	15644
x"00",	-- Hex Addr	3D1D	15645
x"00",	-- Hex Addr	3D1E	15646
x"00",	-- Hex Addr	3D1F	15647
x"00",	-- Hex Addr	3D20	15648
x"00",	-- Hex Addr	3D21	15649
x"00",	-- Hex Addr	3D22	15650
x"00",	-- Hex Addr	3D23	15651
x"00",	-- Hex Addr	3D24	15652
x"00",	-- Hex Addr	3D25	15653
x"00",	-- Hex Addr	3D26	15654
x"00",	-- Hex Addr	3D27	15655
x"00",	-- Hex Addr	3D28	15656
x"00",	-- Hex Addr	3D29	15657
x"00",	-- Hex Addr	3D2A	15658
x"00",	-- Hex Addr	3D2B	15659
x"00",	-- Hex Addr	3D2C	15660
x"00",	-- Hex Addr	3D2D	15661
x"00",	-- Hex Addr	3D2E	15662
x"00",	-- Hex Addr	3D2F	15663
x"00",	-- Hex Addr	3D30	15664
x"00",	-- Hex Addr	3D31	15665
x"00",	-- Hex Addr	3D32	15666
x"00",	-- Hex Addr	3D33	15667
x"00",	-- Hex Addr	3D34	15668
x"00",	-- Hex Addr	3D35	15669
x"00",	-- Hex Addr	3D36	15670
x"00",	-- Hex Addr	3D37	15671
x"00",	-- Hex Addr	3D38	15672
x"00",	-- Hex Addr	3D39	15673
x"00",	-- Hex Addr	3D3A	15674
x"00",	-- Hex Addr	3D3B	15675
x"00",	-- Hex Addr	3D3C	15676
x"00",	-- Hex Addr	3D3D	15677
x"00",	-- Hex Addr	3D3E	15678
x"00",	-- Hex Addr	3D3F	15679
x"00",	-- Hex Addr	3D40	15680
x"00",	-- Hex Addr	3D41	15681
x"00",	-- Hex Addr	3D42	15682
x"00",	-- Hex Addr	3D43	15683
x"00",	-- Hex Addr	3D44	15684
x"00",	-- Hex Addr	3D45	15685
x"00",	-- Hex Addr	3D46	15686
x"00",	-- Hex Addr	3D47	15687
x"00",	-- Hex Addr	3D48	15688
x"00",	-- Hex Addr	3D49	15689
x"00",	-- Hex Addr	3D4A	15690
x"00",	-- Hex Addr	3D4B	15691
x"00",	-- Hex Addr	3D4C	15692
x"00",	-- Hex Addr	3D4D	15693
x"00",	-- Hex Addr	3D4E	15694
x"00",	-- Hex Addr	3D4F	15695
x"00",	-- Hex Addr	3D50	15696
x"00",	-- Hex Addr	3D51	15697
x"00",	-- Hex Addr	3D52	15698
x"00",	-- Hex Addr	3D53	15699
x"00",	-- Hex Addr	3D54	15700
x"00",	-- Hex Addr	3D55	15701
x"00",	-- Hex Addr	3D56	15702
x"00",	-- Hex Addr	3D57	15703
x"00",	-- Hex Addr	3D58	15704
x"00",	-- Hex Addr	3D59	15705
x"00",	-- Hex Addr	3D5A	15706
x"00",	-- Hex Addr	3D5B	15707
x"00",	-- Hex Addr	3D5C	15708
x"00",	-- Hex Addr	3D5D	15709
x"00",	-- Hex Addr	3D5E	15710
x"00",	-- Hex Addr	3D5F	15711
x"00",	-- Hex Addr	3D60	15712
x"00",	-- Hex Addr	3D61	15713
x"00",	-- Hex Addr	3D62	15714
x"00",	-- Hex Addr	3D63	15715
x"00",	-- Hex Addr	3D64	15716
x"00",	-- Hex Addr	3D65	15717
x"00",	-- Hex Addr	3D66	15718
x"00",	-- Hex Addr	3D67	15719
x"00",	-- Hex Addr	3D68	15720
x"00",	-- Hex Addr	3D69	15721
x"00",	-- Hex Addr	3D6A	15722
x"00",	-- Hex Addr	3D6B	15723
x"00",	-- Hex Addr	3D6C	15724
x"00",	-- Hex Addr	3D6D	15725
x"00",	-- Hex Addr	3D6E	15726
x"00",	-- Hex Addr	3D6F	15727
x"00",	-- Hex Addr	3D70	15728
x"00",	-- Hex Addr	3D71	15729
x"00",	-- Hex Addr	3D72	15730
x"00",	-- Hex Addr	3D73	15731
x"00",	-- Hex Addr	3D74	15732
x"00",	-- Hex Addr	3D75	15733
x"00",	-- Hex Addr	3D76	15734
x"00",	-- Hex Addr	3D77	15735
x"00",	-- Hex Addr	3D78	15736
x"00",	-- Hex Addr	3D79	15737
x"00",	-- Hex Addr	3D7A	15738
x"00",	-- Hex Addr	3D7B	15739
x"00",	-- Hex Addr	3D7C	15740
x"00",	-- Hex Addr	3D7D	15741
x"00",	-- Hex Addr	3D7E	15742
x"00",	-- Hex Addr	3D7F	15743
x"00",	-- Hex Addr	3D80	15744
x"00",	-- Hex Addr	3D81	15745
x"00",	-- Hex Addr	3D82	15746
x"00",	-- Hex Addr	3D83	15747
x"00",	-- Hex Addr	3D84	15748
x"00",	-- Hex Addr	3D85	15749
x"00",	-- Hex Addr	3D86	15750
x"00",	-- Hex Addr	3D87	15751
x"00",	-- Hex Addr	3D88	15752
x"00",	-- Hex Addr	3D89	15753
x"00",	-- Hex Addr	3D8A	15754
x"00",	-- Hex Addr	3D8B	15755
x"00",	-- Hex Addr	3D8C	15756
x"00",	-- Hex Addr	3D8D	15757
x"00",	-- Hex Addr	3D8E	15758
x"00",	-- Hex Addr	3D8F	15759
x"00",	-- Hex Addr	3D90	15760
x"00",	-- Hex Addr	3D91	15761
x"00",	-- Hex Addr	3D92	15762
x"00",	-- Hex Addr	3D93	15763
x"00",	-- Hex Addr	3D94	15764
x"00",	-- Hex Addr	3D95	15765
x"00",	-- Hex Addr	3D96	15766
x"00",	-- Hex Addr	3D97	15767
x"00",	-- Hex Addr	3D98	15768
x"00",	-- Hex Addr	3D99	15769
x"00",	-- Hex Addr	3D9A	15770
x"00",	-- Hex Addr	3D9B	15771
x"00",	-- Hex Addr	3D9C	15772
x"00",	-- Hex Addr	3D9D	15773
x"00",	-- Hex Addr	3D9E	15774
x"00",	-- Hex Addr	3D9F	15775
x"00",	-- Hex Addr	3DA0	15776
x"00",	-- Hex Addr	3DA1	15777
x"00",	-- Hex Addr	3DA2	15778
x"00",	-- Hex Addr	3DA3	15779
x"00",	-- Hex Addr	3DA4	15780
x"00",	-- Hex Addr	3DA5	15781
x"00",	-- Hex Addr	3DA6	15782
x"00",	-- Hex Addr	3DA7	15783
x"00",	-- Hex Addr	3DA8	15784
x"00",	-- Hex Addr	3DA9	15785
x"00",	-- Hex Addr	3DAA	15786
x"00",	-- Hex Addr	3DAB	15787
x"00",	-- Hex Addr	3DAC	15788
x"00",	-- Hex Addr	3DAD	15789
x"00",	-- Hex Addr	3DAE	15790
x"00",	-- Hex Addr	3DAF	15791
x"00",	-- Hex Addr	3DB0	15792
x"00",	-- Hex Addr	3DB1	15793
x"00",	-- Hex Addr	3DB2	15794
x"00",	-- Hex Addr	3DB3	15795
x"00",	-- Hex Addr	3DB4	15796
x"00",	-- Hex Addr	3DB5	15797
x"00",	-- Hex Addr	3DB6	15798
x"00",	-- Hex Addr	3DB7	15799
x"00",	-- Hex Addr	3DB8	15800
x"00",	-- Hex Addr	3DB9	15801
x"00",	-- Hex Addr	3DBA	15802
x"00",	-- Hex Addr	3DBB	15803
x"00",	-- Hex Addr	3DBC	15804
x"00",	-- Hex Addr	3DBD	15805
x"00",	-- Hex Addr	3DBE	15806
x"00",	-- Hex Addr	3DBF	15807
x"00",	-- Hex Addr	3DC0	15808
x"00",	-- Hex Addr	3DC1	15809
x"00",	-- Hex Addr	3DC2	15810
x"00",	-- Hex Addr	3DC3	15811
x"00",	-- Hex Addr	3DC4	15812
x"00",	-- Hex Addr	3DC5	15813
x"00",	-- Hex Addr	3DC6	15814
x"00",	-- Hex Addr	3DC7	15815
x"00",	-- Hex Addr	3DC8	15816
x"00",	-- Hex Addr	3DC9	15817
x"00",	-- Hex Addr	3DCA	15818
x"00",	-- Hex Addr	3DCB	15819
x"00",	-- Hex Addr	3DCC	15820
x"00",	-- Hex Addr	3DCD	15821
x"00",	-- Hex Addr	3DCE	15822
x"00",	-- Hex Addr	3DCF	15823
x"00",	-- Hex Addr	3DD0	15824
x"00",	-- Hex Addr	3DD1	15825
x"00",	-- Hex Addr	3DD2	15826
x"00",	-- Hex Addr	3DD3	15827
x"00",	-- Hex Addr	3DD4	15828
x"00",	-- Hex Addr	3DD5	15829
x"00",	-- Hex Addr	3DD6	15830
x"00",	-- Hex Addr	3DD7	15831
x"00",	-- Hex Addr	3DD8	15832
x"00",	-- Hex Addr	3DD9	15833
x"00",	-- Hex Addr	3DDA	15834
x"00",	-- Hex Addr	3DDB	15835
x"00",	-- Hex Addr	3DDC	15836
x"00",	-- Hex Addr	3DDD	15837
x"00",	-- Hex Addr	3DDE	15838
x"00",	-- Hex Addr	3DDF	15839
x"00",	-- Hex Addr	3DE0	15840
x"00",	-- Hex Addr	3DE1	15841
x"00",	-- Hex Addr	3DE2	15842
x"00",	-- Hex Addr	3DE3	15843
x"00",	-- Hex Addr	3DE4	15844
x"00",	-- Hex Addr	3DE5	15845
x"00",	-- Hex Addr	3DE6	15846
x"00",	-- Hex Addr	3DE7	15847
x"00",	-- Hex Addr	3DE8	15848
x"00",	-- Hex Addr	3DE9	15849
x"00",	-- Hex Addr	3DEA	15850
x"00",	-- Hex Addr	3DEB	15851
x"00",	-- Hex Addr	3DEC	15852
x"00",	-- Hex Addr	3DED	15853
x"00",	-- Hex Addr	3DEE	15854
x"00",	-- Hex Addr	3DEF	15855
x"00",	-- Hex Addr	3DF0	15856
x"00",	-- Hex Addr	3DF1	15857
x"00",	-- Hex Addr	3DF2	15858
x"00",	-- Hex Addr	3DF3	15859
x"00",	-- Hex Addr	3DF4	15860
x"00",	-- Hex Addr	3DF5	15861
x"00",	-- Hex Addr	3DF6	15862
x"00",	-- Hex Addr	3DF7	15863
x"00",	-- Hex Addr	3DF8	15864
x"00",	-- Hex Addr	3DF9	15865
x"00",	-- Hex Addr	3DFA	15866
x"00",	-- Hex Addr	3DFB	15867
x"00",	-- Hex Addr	3DFC	15868
x"00",	-- Hex Addr	3DFD	15869
x"00",	-- Hex Addr	3DFE	15870
x"00",	-- Hex Addr	3DFF	15871
x"00",	-- Hex Addr	3E00	15872
x"00",	-- Hex Addr	3E01	15873
x"00",	-- Hex Addr	3E02	15874
x"00",	-- Hex Addr	3E03	15875
x"00",	-- Hex Addr	3E04	15876
x"00",	-- Hex Addr	3E05	15877
x"00",	-- Hex Addr	3E06	15878
x"00",	-- Hex Addr	3E07	15879
x"00",	-- Hex Addr	3E08	15880
x"00",	-- Hex Addr	3E09	15881
x"00",	-- Hex Addr	3E0A	15882
x"00",	-- Hex Addr	3E0B	15883
x"00",	-- Hex Addr	3E0C	15884
x"00",	-- Hex Addr	3E0D	15885
x"00",	-- Hex Addr	3E0E	15886
x"00",	-- Hex Addr	3E0F	15887
x"00",	-- Hex Addr	3E10	15888
x"00",	-- Hex Addr	3E11	15889
x"00",	-- Hex Addr	3E12	15890
x"00",	-- Hex Addr	3E13	15891
x"00",	-- Hex Addr	3E14	15892
x"00",	-- Hex Addr	3E15	15893
x"00",	-- Hex Addr	3E16	15894
x"00",	-- Hex Addr	3E17	15895
x"00",	-- Hex Addr	3E18	15896
x"00",	-- Hex Addr	3E19	15897
x"00",	-- Hex Addr	3E1A	15898
x"00",	-- Hex Addr	3E1B	15899
x"00",	-- Hex Addr	3E1C	15900
x"00",	-- Hex Addr	3E1D	15901
x"00",	-- Hex Addr	3E1E	15902
x"00",	-- Hex Addr	3E1F	15903
x"00",	-- Hex Addr	3E20	15904
x"00",	-- Hex Addr	3E21	15905
x"00",	-- Hex Addr	3E22	15906
x"00",	-- Hex Addr	3E23	15907
x"00",	-- Hex Addr	3E24	15908
x"00",	-- Hex Addr	3E25	15909
x"00",	-- Hex Addr	3E26	15910
x"00",	-- Hex Addr	3E27	15911
x"00",	-- Hex Addr	3E28	15912
x"00",	-- Hex Addr	3E29	15913
x"00",	-- Hex Addr	3E2A	15914
x"00",	-- Hex Addr	3E2B	15915
x"00",	-- Hex Addr	3E2C	15916
x"00",	-- Hex Addr	3E2D	15917
x"00",	-- Hex Addr	3E2E	15918
x"00",	-- Hex Addr	3E2F	15919
x"00",	-- Hex Addr	3E30	15920
x"00",	-- Hex Addr	3E31	15921
x"00",	-- Hex Addr	3E32	15922
x"00",	-- Hex Addr	3E33	15923
x"00",	-- Hex Addr	3E34	15924
x"00",	-- Hex Addr	3E35	15925
x"00",	-- Hex Addr	3E36	15926
x"00",	-- Hex Addr	3E37	15927
x"00",	-- Hex Addr	3E38	15928
x"00",	-- Hex Addr	3E39	15929
x"00",	-- Hex Addr	3E3A	15930
x"00",	-- Hex Addr	3E3B	15931
x"00",	-- Hex Addr	3E3C	15932
x"00",	-- Hex Addr	3E3D	15933
x"00",	-- Hex Addr	3E3E	15934
x"00",	-- Hex Addr	3E3F	15935
x"00",	-- Hex Addr	3E40	15936
x"00",	-- Hex Addr	3E41	15937
x"00",	-- Hex Addr	3E42	15938
x"00",	-- Hex Addr	3E43	15939
x"00",	-- Hex Addr	3E44	15940
x"00",	-- Hex Addr	3E45	15941
x"00",	-- Hex Addr	3E46	15942
x"00",	-- Hex Addr	3E47	15943
x"00",	-- Hex Addr	3E48	15944
x"00",	-- Hex Addr	3E49	15945
x"00",	-- Hex Addr	3E4A	15946
x"00",	-- Hex Addr	3E4B	15947
x"00",	-- Hex Addr	3E4C	15948
x"00",	-- Hex Addr	3E4D	15949
x"00",	-- Hex Addr	3E4E	15950
x"00",	-- Hex Addr	3E4F	15951
x"00",	-- Hex Addr	3E50	15952
x"00",	-- Hex Addr	3E51	15953
x"00",	-- Hex Addr	3E52	15954
x"00",	-- Hex Addr	3E53	15955
x"00",	-- Hex Addr	3E54	15956
x"00",	-- Hex Addr	3E55	15957
x"00",	-- Hex Addr	3E56	15958
x"00",	-- Hex Addr	3E57	15959
x"00",	-- Hex Addr	3E58	15960
x"00",	-- Hex Addr	3E59	15961
x"00",	-- Hex Addr	3E5A	15962
x"00",	-- Hex Addr	3E5B	15963
x"00",	-- Hex Addr	3E5C	15964
x"00",	-- Hex Addr	3E5D	15965
x"00",	-- Hex Addr	3E5E	15966
x"00",	-- Hex Addr	3E5F	15967
x"00",	-- Hex Addr	3E60	15968
x"00",	-- Hex Addr	3E61	15969
x"00",	-- Hex Addr	3E62	15970
x"00",	-- Hex Addr	3E63	15971
x"00",	-- Hex Addr	3E64	15972
x"00",	-- Hex Addr	3E65	15973
x"00",	-- Hex Addr	3E66	15974
x"00",	-- Hex Addr	3E67	15975
x"00",	-- Hex Addr	3E68	15976
x"00",	-- Hex Addr	3E69	15977
x"00",	-- Hex Addr	3E6A	15978
x"00",	-- Hex Addr	3E6B	15979
x"00",	-- Hex Addr	3E6C	15980
x"00",	-- Hex Addr	3E6D	15981
x"00",	-- Hex Addr	3E6E	15982
x"00",	-- Hex Addr	3E6F	15983
x"01",	-- Hex Addr	3E70	15984
x"07",	-- Hex Addr	3E71	15985
x"00",	-- Hex Addr	3E72	15986
x"01",	-- Hex Addr	3E73	15987
x"03",	-- Hex Addr	3E74	15988
x"03",	-- Hex Addr	3E75	15989
x"04",	-- Hex Addr	3E76	15990
x"02",	-- Hex Addr	3E77	15991
x"00",	-- Hex Addr	3E78	15992
x"05",	-- Hex Addr	3E79	15993
x"00",	-- Hex Addr	3E7A	15994
x"00",	-- Hex Addr	3E7B	15995
x"00",	-- Hex Addr	3E7C	15996
x"00",	-- Hex Addr	3E7D	15997
x"00",	-- Hex Addr	3E7E	15998
x"00",	-- Hex Addr	3E7F	15999
x"00",	-- Hex Addr	3E80	16000
x"00",	-- Hex Addr	3E81	16001
x"00",	-- Hex Addr	3E82	16002
x"00",	-- Hex Addr	3E83	16003
x"00",	-- Hex Addr	3E84	16004
x"00",	-- Hex Addr	3E85	16005
x"00",	-- Hex Addr	3E86	16006
x"00",	-- Hex Addr	3E87	16007
x"00",	-- Hex Addr	3E88	16008
x"00",	-- Hex Addr	3E89	16009
x"00",	-- Hex Addr	3E8A	16010
x"00",	-- Hex Addr	3E8B	16011
x"00",	-- Hex Addr	3E8C	16012
x"00",	-- Hex Addr	3E8D	16013
x"00",	-- Hex Addr	3E8E	16014
x"00",	-- Hex Addr	3E8F	16015
x"00",	-- Hex Addr	3E90	16016
x"00",	-- Hex Addr	3E91	16017
x"00",	-- Hex Addr	3E92	16018
x"00",	-- Hex Addr	3E93	16019
x"00",	-- Hex Addr	3E94	16020
x"00",	-- Hex Addr	3E95	16021
x"00",	-- Hex Addr	3E96	16022
x"00",	-- Hex Addr	3E97	16023
x"00",	-- Hex Addr	3E98	16024
x"00",	-- Hex Addr	3E99	16025
x"00",	-- Hex Addr	3E9A	16026
x"00",	-- Hex Addr	3E9B	16027
x"00",	-- Hex Addr	3E9C	16028
x"00",	-- Hex Addr	3E9D	16029
x"00",	-- Hex Addr	3E9E	16030
x"00",	-- Hex Addr	3E9F	16031
x"00",	-- Hex Addr	3EA0	16032
x"00",	-- Hex Addr	3EA1	16033
x"00",	-- Hex Addr	3EA2	16034
x"00",	-- Hex Addr	3EA3	16035
x"00",	-- Hex Addr	3EA4	16036
x"00",	-- Hex Addr	3EA5	16037
x"00",	-- Hex Addr	3EA6	16038
x"00",	-- Hex Addr	3EA7	16039
x"00",	-- Hex Addr	3EA8	16040
x"00",	-- Hex Addr	3EA9	16041
x"00",	-- Hex Addr	3EAA	16042
x"00",	-- Hex Addr	3EAB	16043
x"00",	-- Hex Addr	3EAC	16044
x"00",	-- Hex Addr	3EAD	16045
x"00",	-- Hex Addr	3EAE	16046
x"00",	-- Hex Addr	3EAF	16047
x"00",	-- Hex Addr	3EB0	16048
x"00",	-- Hex Addr	3EB1	16049
x"00",	-- Hex Addr	3EB2	16050
x"00",	-- Hex Addr	3EB3	16051
x"00",	-- Hex Addr	3EB4	16052
x"00",	-- Hex Addr	3EB5	16053
x"00",	-- Hex Addr	3EB6	16054
x"00",	-- Hex Addr	3EB7	16055
x"00",	-- Hex Addr	3EB8	16056
x"00",	-- Hex Addr	3EB9	16057
x"00",	-- Hex Addr	3EBA	16058
x"00",	-- Hex Addr	3EBB	16059
x"00",	-- Hex Addr	3EBC	16060
x"00",	-- Hex Addr	3EBD	16061
x"00",	-- Hex Addr	3EBE	16062
x"00",	-- Hex Addr	3EBF	16063
x"00",	-- Hex Addr	3EC0	16064
x"00",	-- Hex Addr	3EC1	16065
x"00",	-- Hex Addr	3EC2	16066
x"00",	-- Hex Addr	3EC3	16067
x"00",	-- Hex Addr	3EC4	16068
x"00",	-- Hex Addr	3EC5	16069
x"00",	-- Hex Addr	3EC6	16070
x"00",	-- Hex Addr	3EC7	16071
x"00",	-- Hex Addr	3EC8	16072
x"00",	-- Hex Addr	3EC9	16073
x"00",	-- Hex Addr	3ECA	16074
x"00",	-- Hex Addr	3ECB	16075
x"00",	-- Hex Addr	3ECC	16076
x"00",	-- Hex Addr	3ECD	16077
x"00",	-- Hex Addr	3ECE	16078
x"00",	-- Hex Addr	3ECF	16079
x"00",	-- Hex Addr	3ED0	16080
x"00",	-- Hex Addr	3ED1	16081
x"00",	-- Hex Addr	3ED2	16082
x"00",	-- Hex Addr	3ED3	16083
x"00",	-- Hex Addr	3ED4	16084
x"00",	-- Hex Addr	3ED5	16085
x"00",	-- Hex Addr	3ED6	16086
x"00",	-- Hex Addr	3ED7	16087
x"00",	-- Hex Addr	3ED8	16088
x"00",	-- Hex Addr	3ED9	16089
x"00",	-- Hex Addr	3EDA	16090
x"00",	-- Hex Addr	3EDB	16091
x"00",	-- Hex Addr	3EDC	16092
x"00",	-- Hex Addr	3EDD	16093
x"00",	-- Hex Addr	3EDE	16094
x"00",	-- Hex Addr	3EDF	16095
x"00",	-- Hex Addr	3EE0	16096
x"00",	-- Hex Addr	3EE1	16097
x"00",	-- Hex Addr	3EE2	16098
x"00",	-- Hex Addr	3EE3	16099
x"00",	-- Hex Addr	3EE4	16100
x"00",	-- Hex Addr	3EE5	16101
x"00",	-- Hex Addr	3EE6	16102
x"00",	-- Hex Addr	3EE7	16103
x"00",	-- Hex Addr	3EE8	16104
x"00",	-- Hex Addr	3EE9	16105
x"00",	-- Hex Addr	3EEA	16106
x"00",	-- Hex Addr	3EEB	16107
x"00",	-- Hex Addr	3EEC	16108
x"00",	-- Hex Addr	3EED	16109
x"00",	-- Hex Addr	3EEE	16110
x"00",	-- Hex Addr	3EEF	16111
x"00",	-- Hex Addr	3EF0	16112
x"00",	-- Hex Addr	3EF1	16113
x"00",	-- Hex Addr	3EF2	16114
x"00",	-- Hex Addr	3EF3	16115
x"00",	-- Hex Addr	3EF4	16116
x"00",	-- Hex Addr	3EF5	16117
x"00",	-- Hex Addr	3EF6	16118
x"00",	-- Hex Addr	3EF7	16119
x"00",	-- Hex Addr	3EF8	16120
x"00",	-- Hex Addr	3EF9	16121
x"00",	-- Hex Addr	3EFA	16122
x"00",	-- Hex Addr	3EFB	16123
x"00",	-- Hex Addr	3EFC	16124
x"00",	-- Hex Addr	3EFD	16125
x"00",	-- Hex Addr	3EFE	16126
x"00",	-- Hex Addr	3EFF	16127
x"00",	-- Hex Addr	3F00	16128
x"00",	-- Hex Addr	3F01	16129
x"00",	-- Hex Addr	3F02	16130
x"00",	-- Hex Addr	3F03	16131
x"00",	-- Hex Addr	3F04	16132
x"00",	-- Hex Addr	3F05	16133
x"00",	-- Hex Addr	3F06	16134
x"00",	-- Hex Addr	3F07	16135
x"00",	-- Hex Addr	3F08	16136
x"00",	-- Hex Addr	3F09	16137
x"00",	-- Hex Addr	3F0A	16138
x"00",	-- Hex Addr	3F0B	16139
x"00",	-- Hex Addr	3F0C	16140
x"00",	-- Hex Addr	3F0D	16141
x"00",	-- Hex Addr	3F0E	16142
x"00",	-- Hex Addr	3F0F	16143
x"00",	-- Hex Addr	3F10	16144
x"00",	-- Hex Addr	3F11	16145
x"00",	-- Hex Addr	3F12	16146
x"00",	-- Hex Addr	3F13	16147
x"00",	-- Hex Addr	3F14	16148
x"00",	-- Hex Addr	3F15	16149
x"00",	-- Hex Addr	3F16	16150
x"00",	-- Hex Addr	3F17	16151
x"00",	-- Hex Addr	3F18	16152
x"00",	-- Hex Addr	3F19	16153
x"00",	-- Hex Addr	3F1A	16154
x"00",	-- Hex Addr	3F1B	16155
x"00",	-- Hex Addr	3F1C	16156
x"00",	-- Hex Addr	3F1D	16157
x"00",	-- Hex Addr	3F1E	16158
x"00",	-- Hex Addr	3F1F	16159
x"00",	-- Hex Addr	3F20	16160
x"00",	-- Hex Addr	3F21	16161
x"00",	-- Hex Addr	3F22	16162
x"00",	-- Hex Addr	3F23	16163
x"00",	-- Hex Addr	3F24	16164
x"00",	-- Hex Addr	3F25	16165
x"00",	-- Hex Addr	3F26	16166
x"00",	-- Hex Addr	3F27	16167
x"00",	-- Hex Addr	3F28	16168
x"00",	-- Hex Addr	3F29	16169
x"00",	-- Hex Addr	3F2A	16170
x"00",	-- Hex Addr	3F2B	16171
x"00",	-- Hex Addr	3F2C	16172
x"00",	-- Hex Addr	3F2D	16173
x"00",	-- Hex Addr	3F2E	16174
x"00",	-- Hex Addr	3F2F	16175
x"00",	-- Hex Addr	3F30	16176
x"00",	-- Hex Addr	3F31	16177
x"00",	-- Hex Addr	3F32	16178
x"00",	-- Hex Addr	3F33	16179
x"00",	-- Hex Addr	3F34	16180
x"00",	-- Hex Addr	3F35	16181
x"00",	-- Hex Addr	3F36	16182
x"00",	-- Hex Addr	3F37	16183
x"00",	-- Hex Addr	3F38	16184
x"00",	-- Hex Addr	3F39	16185
x"00",	-- Hex Addr	3F3A	16186
x"00",	-- Hex Addr	3F3B	16187
x"00",	-- Hex Addr	3F3C	16188
x"00",	-- Hex Addr	3F3D	16189
x"00",	-- Hex Addr	3F3E	16190
x"00",	-- Hex Addr	3F3F	16191
x"00",	-- Hex Addr	3F40	16192
x"00",	-- Hex Addr	3F41	16193
x"00",	-- Hex Addr	3F42	16194
x"00",	-- Hex Addr	3F43	16195
x"00",	-- Hex Addr	3F44	16196
x"00",	-- Hex Addr	3F45	16197
x"00",	-- Hex Addr	3F46	16198
x"00",	-- Hex Addr	3F47	16199
x"00",	-- Hex Addr	3F48	16200
x"00",	-- Hex Addr	3F49	16201
x"00",	-- Hex Addr	3F4A	16202
x"00",	-- Hex Addr	3F4B	16203
x"00",	-- Hex Addr	3F4C	16204
x"00",	-- Hex Addr	3F4D	16205
x"00",	-- Hex Addr	3F4E	16206
x"00",	-- Hex Addr	3F4F	16207
x"00",	-- Hex Addr	3F50	16208
x"00",	-- Hex Addr	3F51	16209
x"00",	-- Hex Addr	3F52	16210
x"00",	-- Hex Addr	3F53	16211
x"00",	-- Hex Addr	3F54	16212
x"00",	-- Hex Addr	3F55	16213
x"00",	-- Hex Addr	3F56	16214
x"00",	-- Hex Addr	3F57	16215
x"00",	-- Hex Addr	3F58	16216
x"00",	-- Hex Addr	3F59	16217
x"00",	-- Hex Addr	3F5A	16218
x"00",	-- Hex Addr	3F5B	16219
x"00",	-- Hex Addr	3F5C	16220
x"00",	-- Hex Addr	3F5D	16221
x"00",	-- Hex Addr	3F5E	16222
x"00",	-- Hex Addr	3F5F	16223
x"00",	-- Hex Addr	3F60	16224
x"00",	-- Hex Addr	3F61	16225
x"00",	-- Hex Addr	3F62	16226
x"00",	-- Hex Addr	3F63	16227
x"00",	-- Hex Addr	3F64	16228
x"00",	-- Hex Addr	3F65	16229
x"00",	-- Hex Addr	3F66	16230
x"00",	-- Hex Addr	3F67	16231
x"00",	-- Hex Addr	3F68	16232
x"00",	-- Hex Addr	3F69	16233
x"00",	-- Hex Addr	3F6A	16234
x"00",	-- Hex Addr	3F6B	16235
x"00",	-- Hex Addr	3F6C	16236
x"00",	-- Hex Addr	3F6D	16237
x"00",	-- Hex Addr	3F6E	16238
x"00",	-- Hex Addr	3F6F	16239
x"00",	-- Hex Addr	3F70	16240
x"00",	-- Hex Addr	3F71	16241
x"00",	-- Hex Addr	3F72	16242
x"00",	-- Hex Addr	3F73	16243
x"00",	-- Hex Addr	3F74	16244
x"00",	-- Hex Addr	3F75	16245
x"00",	-- Hex Addr	3F76	16246
x"00",	-- Hex Addr	3F77	16247
x"00",	-- Hex Addr	3F78	16248
x"00",	-- Hex Addr	3F79	16249
x"00",	-- Hex Addr	3F7A	16250
x"00",	-- Hex Addr	3F7B	16251
x"00",	-- Hex Addr	3F7C	16252
x"00",	-- Hex Addr	3F7D	16253
x"00",	-- Hex Addr	3F7E	16254
x"00",	-- Hex Addr	3F7F	16255
x"00",	-- Hex Addr	3F80	16256
x"00",	-- Hex Addr	3F81	16257
x"00",	-- Hex Addr	3F82	16258
x"00",	-- Hex Addr	3F83	16259
x"00",	-- Hex Addr	3F84	16260
x"00",	-- Hex Addr	3F85	16261
x"00",	-- Hex Addr	3F86	16262
x"00",	-- Hex Addr	3F87	16263
x"00",	-- Hex Addr	3F88	16264
x"00",	-- Hex Addr	3F89	16265
x"00",	-- Hex Addr	3F8A	16266
x"00",	-- Hex Addr	3F8B	16267
x"00",	-- Hex Addr	3F8C	16268
x"00",	-- Hex Addr	3F8D	16269
x"00",	-- Hex Addr	3F8E	16270
x"00",	-- Hex Addr	3F8F	16271
x"00",	-- Hex Addr	3F90	16272
x"00",	-- Hex Addr	3F91	16273
x"00",	-- Hex Addr	3F92	16274
x"00",	-- Hex Addr	3F93	16275
x"00",	-- Hex Addr	3F94	16276
x"00",	-- Hex Addr	3F95	16277
x"00",	-- Hex Addr	3F96	16278
x"00",	-- Hex Addr	3F97	16279
x"00",	-- Hex Addr	3F98	16280
x"00",	-- Hex Addr	3F99	16281
x"00",	-- Hex Addr	3F9A	16282
x"00",	-- Hex Addr	3F9B	16283
x"00",	-- Hex Addr	3F9C	16284
x"00",	-- Hex Addr	3F9D	16285
x"00",	-- Hex Addr	3F9E	16286
x"00",	-- Hex Addr	3F9F	16287
x"00",	-- Hex Addr	3FA0	16288
x"00",	-- Hex Addr	3FA1	16289
x"00",	-- Hex Addr	3FA2	16290
x"00",	-- Hex Addr	3FA3	16291
x"00",	-- Hex Addr	3FA4	16292
x"00",	-- Hex Addr	3FA5	16293
x"00",	-- Hex Addr	3FA6	16294
x"00",	-- Hex Addr	3FA7	16295
x"00",	-- Hex Addr	3FA8	16296
x"00",	-- Hex Addr	3FA9	16297
x"00",	-- Hex Addr	3FAA	16298
x"00",	-- Hex Addr	3FAB	16299
x"00",	-- Hex Addr	3FAC	16300
x"00",	-- Hex Addr	3FAD	16301
x"00",	-- Hex Addr	3FAE	16302
x"00",	-- Hex Addr	3FAF	16303
x"00",	-- Hex Addr	3FB0	16304
x"00",	-- Hex Addr	3FB1	16305
x"00",	-- Hex Addr	3FB2	16306
x"00",	-- Hex Addr	3FB3	16307
x"00",	-- Hex Addr	3FB4	16308
x"00",	-- Hex Addr	3FB5	16309
x"00",	-- Hex Addr	3FB6	16310
x"00",	-- Hex Addr	3FB7	16311
x"00",	-- Hex Addr	3FB8	16312
x"00",	-- Hex Addr	3FB9	16313
x"00",	-- Hex Addr	3FBA	16314
x"00",	-- Hex Addr	3FBB	16315
x"00",	-- Hex Addr	3FBC	16316
x"00",	-- Hex Addr	3FBD	16317
x"00",	-- Hex Addr	3FBE	16318
x"00",	-- Hex Addr	3FBF	16319
x"00",	-- Hex Addr	3FC0	16320
x"00",	-- Hex Addr	3FC1	16321
x"00",	-- Hex Addr	3FC2	16322
x"00",	-- Hex Addr	3FC3	16323
x"00",	-- Hex Addr	3FC4	16324
x"00",	-- Hex Addr	3FC5	16325
x"00",	-- Hex Addr	3FC6	16326
x"00",	-- Hex Addr	3FC7	16327
x"00",	-- Hex Addr	3FC8	16328
x"00",	-- Hex Addr	3FC9	16329
x"00",	-- Hex Addr	3FCA	16330
x"00",	-- Hex Addr	3FCB	16331
x"00",	-- Hex Addr	3FCC	16332
x"00",	-- Hex Addr	3FCD	16333
x"00",	-- Hex Addr	3FCE	16334
x"00",	-- Hex Addr	3FCF	16335
x"00",	-- Hex Addr	3FD0	16336
x"00",	-- Hex Addr	3FD1	16337
x"00",	-- Hex Addr	3FD2	16338
x"00",	-- Hex Addr	3FD3	16339
x"00",	-- Hex Addr	3FD4	16340
x"00",	-- Hex Addr	3FD5	16341
x"00",	-- Hex Addr	3FD6	16342
x"00",	-- Hex Addr	3FD7	16343
x"00",	-- Hex Addr	3FD8	16344
x"00",	-- Hex Addr	3FD9	16345
x"00",	-- Hex Addr	3FDA	16346
x"00",	-- Hex Addr	3FDB	16347
x"00",	-- Hex Addr	3FDC	16348
x"00",	-- Hex Addr	3FDD	16349
x"00",	-- Hex Addr	3FDE	16350
x"00",	-- Hex Addr	3FDF	16351
x"00",	-- Hex Addr	3FE0	16352
x"00",	-- Hex Addr	3FE1	16353
x"00",	-- Hex Addr	3FE2	16354
x"00",	-- Hex Addr	3FE3	16355
x"00",	-- Hex Addr	3FE4	16356
x"00",	-- Hex Addr	3FE5	16357
x"00",	-- Hex Addr	3FE6	16358
x"00",	-- Hex Addr	3FE7	16359
x"00",	-- Hex Addr	3FE8	16360
x"00",	-- Hex Addr	3FE9	16361
x"00",	-- Hex Addr	3FEA	16362
x"00",	-- Hex Addr	3FEB	16363
x"00",	-- Hex Addr	3FEC	16364
x"00",	-- Hex Addr	3FED	16365
x"00",	-- Hex Addr	3FEE	16366
x"00",	-- Hex Addr	3FEF	16367
x"00",	-- Hex Addr	3FF0	16368
x"00",	-- Hex Addr	3FF1	16369
x"00",	-- Hex Addr	3FF2	16370
x"00",	-- Hex Addr	3FF3	16371
x"00",	-- Hex Addr	3FF4	16372
x"00",	-- Hex Addr	3FF5	16373
x"00",	-- Hex Addr	3FF6	16374
x"00",	-- Hex Addr	3FF7	16375
x"00",	-- Hex Addr	3FF8	16376
x"00",	-- Hex Addr	3FF9	16377
x"00",	-- Hex Addr	3FFA	16378
x"00",	-- Hex Addr	3FFB	16379
x"00",	-- Hex Addr	3FFC	16380
x"00",	-- Hex Addr	3FFD	16381
x"00",	-- Hex Addr	3FFE	16382
x"00",	-- Hex Addr	3FFF	16383
x"00",	-- Hex Addr	4000	16384
x"00",	-- Hex Addr	4001	16385
x"00",	-- Hex Addr	4002	16386
x"00",	-- Hex Addr	4003	16387
x"00",	-- Hex Addr	4004	16388
x"00",	-- Hex Addr	4005	16389
x"00",	-- Hex Addr	4006	16390
x"00",	-- Hex Addr	4007	16391
x"00",	-- Hex Addr	4008	16392
x"00",	-- Hex Addr	4009	16393
x"00",	-- Hex Addr	400A	16394
x"00",	-- Hex Addr	400B	16395
x"00",	-- Hex Addr	400C	16396
x"00",	-- Hex Addr	400D	16397
x"00",	-- Hex Addr	400E	16398
x"00",	-- Hex Addr	400F	16399
x"00",	-- Hex Addr	4010	16400
x"00",	-- Hex Addr	4011	16401
x"00",	-- Hex Addr	4012	16402
x"00",	-- Hex Addr	4013	16403
x"00",	-- Hex Addr	4014	16404
x"00",	-- Hex Addr	4015	16405
x"00",	-- Hex Addr	4016	16406
x"00",	-- Hex Addr	4017	16407
x"00",	-- Hex Addr	4018	16408
x"00",	-- Hex Addr	4019	16409
x"00",	-- Hex Addr	401A	16410
x"00",	-- Hex Addr	401B	16411
x"00",	-- Hex Addr	401C	16412
x"00",	-- Hex Addr	401D	16413
x"00",	-- Hex Addr	401E	16414
x"00",	-- Hex Addr	401F	16415
x"00",	-- Hex Addr	4020	16416
x"00",	-- Hex Addr	4021	16417
x"00",	-- Hex Addr	4022	16418
x"00",	-- Hex Addr	4023	16419
x"00",	-- Hex Addr	4024	16420
x"00",	-- Hex Addr	4025	16421
x"00",	-- Hex Addr	4026	16422
x"00",	-- Hex Addr	4027	16423
x"00",	-- Hex Addr	4028	16424
x"00",	-- Hex Addr	4029	16425
x"00",	-- Hex Addr	402A	16426
x"00",	-- Hex Addr	402B	16427
x"00",	-- Hex Addr	402C	16428
x"00",	-- Hex Addr	402D	16429
x"00",	-- Hex Addr	402E	16430
x"00",	-- Hex Addr	402F	16431
x"00",	-- Hex Addr	4030	16432
x"00",	-- Hex Addr	4031	16433
x"00",	-- Hex Addr	4032	16434
x"00",	-- Hex Addr	4033	16435
x"00",	-- Hex Addr	4034	16436
x"00",	-- Hex Addr	4035	16437
x"00",	-- Hex Addr	4036	16438
x"00",	-- Hex Addr	4037	16439
x"00",	-- Hex Addr	4038	16440
x"00",	-- Hex Addr	4039	16441
x"00",	-- Hex Addr	403A	16442
x"00",	-- Hex Addr	403B	16443
x"00",	-- Hex Addr	403C	16444
x"00",	-- Hex Addr	403D	16445
x"00",	-- Hex Addr	403E	16446
x"00",	-- Hex Addr	403F	16447
x"00",	-- Hex Addr	4040	16448
x"00",	-- Hex Addr	4041	16449
x"00",	-- Hex Addr	4042	16450
x"00",	-- Hex Addr	4043	16451
x"00",	-- Hex Addr	4044	16452
x"00",	-- Hex Addr	4045	16453
x"00",	-- Hex Addr	4046	16454
x"00",	-- Hex Addr	4047	16455
x"00",	-- Hex Addr	4048	16456
x"00",	-- Hex Addr	4049	16457
x"00",	-- Hex Addr	404A	16458
x"00",	-- Hex Addr	404B	16459
x"00",	-- Hex Addr	404C	16460
x"00",	-- Hex Addr	404D	16461
x"00",	-- Hex Addr	404E	16462
x"00",	-- Hex Addr	404F	16463
x"00",	-- Hex Addr	4050	16464
x"00",	-- Hex Addr	4051	16465
x"00",	-- Hex Addr	4052	16466
x"00",	-- Hex Addr	4053	16467
x"00",	-- Hex Addr	4054	16468
x"00",	-- Hex Addr	4055	16469
x"00",	-- Hex Addr	4056	16470
x"00",	-- Hex Addr	4057	16471
x"00",	-- Hex Addr	4058	16472
x"00",	-- Hex Addr	4059	16473
x"00",	-- Hex Addr	405A	16474
x"00",	-- Hex Addr	405B	16475
x"00",	-- Hex Addr	405C	16476
x"00",	-- Hex Addr	405D	16477
x"00",	-- Hex Addr	405E	16478
x"00",	-- Hex Addr	405F	16479
x"00",	-- Hex Addr	4060	16480
x"00",	-- Hex Addr	4061	16481
x"00",	-- Hex Addr	4062	16482
x"00",	-- Hex Addr	4063	16483
x"00",	-- Hex Addr	4064	16484
x"00",	-- Hex Addr	4065	16485
x"00",	-- Hex Addr	4066	16486
x"00",	-- Hex Addr	4067	16487
x"00",	-- Hex Addr	4068	16488
x"00",	-- Hex Addr	4069	16489
x"00",	-- Hex Addr	406A	16490
x"00",	-- Hex Addr	406B	16491
x"00",	-- Hex Addr	406C	16492
x"00",	-- Hex Addr	406D	16493
x"00",	-- Hex Addr	406E	16494
x"00",	-- Hex Addr	406F	16495
x"00",	-- Hex Addr	4070	16496
x"00",	-- Hex Addr	4071	16497
x"00",	-- Hex Addr	4072	16498
x"00",	-- Hex Addr	4073	16499
x"00",	-- Hex Addr	4074	16500
x"00",	-- Hex Addr	4075	16501
x"00",	-- Hex Addr	4076	16502
x"00",	-- Hex Addr	4077	16503
x"00",	-- Hex Addr	4078	16504
x"00",	-- Hex Addr	4079	16505
x"00",	-- Hex Addr	407A	16506
x"00",	-- Hex Addr	407B	16507
x"00",	-- Hex Addr	407C	16508
x"00",	-- Hex Addr	407D	16509
x"00",	-- Hex Addr	407E	16510
x"00",	-- Hex Addr	407F	16511
x"00",	-- Hex Addr	4080	16512
x"00",	-- Hex Addr	4081	16513
x"00",	-- Hex Addr	4082	16514
x"00",	-- Hex Addr	4083	16515
x"00",	-- Hex Addr	4084	16516
x"00",	-- Hex Addr	4085	16517
x"00",	-- Hex Addr	4086	16518
x"00",	-- Hex Addr	4087	16519
x"00",	-- Hex Addr	4088	16520
x"00",	-- Hex Addr	4089	16521
x"00",	-- Hex Addr	408A	16522
x"00",	-- Hex Addr	408B	16523
x"00",	-- Hex Addr	408C	16524
x"00",	-- Hex Addr	408D	16525
x"00",	-- Hex Addr	408E	16526
x"00",	-- Hex Addr	408F	16527
x"00",	-- Hex Addr	4090	16528
x"00",	-- Hex Addr	4091	16529
x"00",	-- Hex Addr	4092	16530
x"00",	-- Hex Addr	4093	16531
x"00",	-- Hex Addr	4094	16532
x"00",	-- Hex Addr	4095	16533
x"00",	-- Hex Addr	4096	16534
x"00",	-- Hex Addr	4097	16535
x"00",	-- Hex Addr	4098	16536
x"00",	-- Hex Addr	4099	16537
x"00",	-- Hex Addr	409A	16538
x"00",	-- Hex Addr	409B	16539
x"00",	-- Hex Addr	409C	16540
x"00",	-- Hex Addr	409D	16541
x"00",	-- Hex Addr	409E	16542
x"00",	-- Hex Addr	409F	16543
x"00",	-- Hex Addr	40A0	16544
x"00",	-- Hex Addr	40A1	16545
x"00",	-- Hex Addr	40A2	16546
x"00",	-- Hex Addr	40A3	16547
x"00",	-- Hex Addr	40A4	16548
x"00",	-- Hex Addr	40A5	16549
x"00",	-- Hex Addr	40A6	16550
x"00",	-- Hex Addr	40A7	16551
x"00",	-- Hex Addr	40A8	16552
x"00",	-- Hex Addr	40A9	16553
x"00",	-- Hex Addr	40AA	16554
x"00",	-- Hex Addr	40AB	16555
x"00",	-- Hex Addr	40AC	16556
x"00",	-- Hex Addr	40AD	16557
x"00",	-- Hex Addr	40AE	16558
x"00",	-- Hex Addr	40AF	16559
x"00",	-- Hex Addr	40B0	16560
x"00",	-- Hex Addr	40B1	16561
x"00",	-- Hex Addr	40B2	16562
x"00",	-- Hex Addr	40B3	16563
x"00",	-- Hex Addr	40B4	16564
x"00",	-- Hex Addr	40B5	16565
x"00",	-- Hex Addr	40B6	16566
x"00",	-- Hex Addr	40B7	16567
x"00",	-- Hex Addr	40B8	16568
x"00",	-- Hex Addr	40B9	16569
x"00",	-- Hex Addr	40BA	16570
x"00",	-- Hex Addr	40BB	16571
x"00",	-- Hex Addr	40BC	16572
x"00",	-- Hex Addr	40BD	16573
x"00",	-- Hex Addr	40BE	16574
x"00",	-- Hex Addr	40BF	16575
x"00",	-- Hex Addr	40C0	16576
x"00",	-- Hex Addr	40C1	16577
x"00",	-- Hex Addr	40C2	16578
x"00",	-- Hex Addr	40C3	16579
x"00",	-- Hex Addr	40C4	16580
x"00",	-- Hex Addr	40C5	16581
x"00",	-- Hex Addr	40C6	16582
x"00",	-- Hex Addr	40C7	16583
x"00",	-- Hex Addr	40C8	16584
x"00",	-- Hex Addr	40C9	16585
x"00",	-- Hex Addr	40CA	16586
x"00",	-- Hex Addr	40CB	16587
x"00",	-- Hex Addr	40CC	16588
x"00",	-- Hex Addr	40CD	16589
x"00",	-- Hex Addr	40CE	16590
x"00",	-- Hex Addr	40CF	16591
x"00",	-- Hex Addr	40D0	16592
x"00",	-- Hex Addr	40D1	16593
x"00",	-- Hex Addr	40D2	16594
x"00",	-- Hex Addr	40D3	16595
x"00",	-- Hex Addr	40D4	16596
x"00",	-- Hex Addr	40D5	16597
x"00",	-- Hex Addr	40D6	16598
x"00",	-- Hex Addr	40D7	16599
x"00",	-- Hex Addr	40D8	16600
x"00",	-- Hex Addr	40D9	16601
x"00",	-- Hex Addr	40DA	16602
x"00",	-- Hex Addr	40DB	16603
x"00",	-- Hex Addr	40DC	16604
x"00",	-- Hex Addr	40DD	16605
x"00",	-- Hex Addr	40DE	16606
x"00",	-- Hex Addr	40DF	16607
x"00",	-- Hex Addr	40E0	16608
x"00",	-- Hex Addr	40E1	16609
x"00",	-- Hex Addr	40E2	16610
x"00",	-- Hex Addr	40E3	16611
x"00",	-- Hex Addr	40E4	16612
x"00",	-- Hex Addr	40E5	16613
x"00",	-- Hex Addr	40E6	16614
x"00",	-- Hex Addr	40E7	16615
x"00",	-- Hex Addr	40E8	16616
x"00",	-- Hex Addr	40E9	16617
x"00",	-- Hex Addr	40EA	16618
x"00",	-- Hex Addr	40EB	16619
x"00",	-- Hex Addr	40EC	16620
x"00",	-- Hex Addr	40ED	16621
x"00",	-- Hex Addr	40EE	16622
x"00",	-- Hex Addr	40EF	16623
x"00",	-- Hex Addr	40F0	16624
x"00",	-- Hex Addr	40F1	16625
x"00",	-- Hex Addr	40F2	16626
x"00",	-- Hex Addr	40F3	16627
x"00",	-- Hex Addr	40F4	16628
x"00",	-- Hex Addr	40F5	16629
x"00",	-- Hex Addr	40F6	16630
x"00",	-- Hex Addr	40F7	16631
x"00",	-- Hex Addr	40F8	16632
x"00",	-- Hex Addr	40F9	16633
x"00",	-- Hex Addr	40FA	16634
x"00",	-- Hex Addr	40FB	16635
x"00",	-- Hex Addr	40FC	16636
x"00",	-- Hex Addr	40FD	16637
x"00",	-- Hex Addr	40FE	16638
x"00",	-- Hex Addr	40FF	16639
x"00",	-- Hex Addr	4100	16640
x"00",	-- Hex Addr	4101	16641
x"00",	-- Hex Addr	4102	16642
x"00",	-- Hex Addr	4103	16643
x"00",	-- Hex Addr	4104	16644
x"00",	-- Hex Addr	4105	16645
x"00",	-- Hex Addr	4106	16646
x"00",	-- Hex Addr	4107	16647
x"00",	-- Hex Addr	4108	16648
x"00",	-- Hex Addr	4109	16649
x"00",	-- Hex Addr	410A	16650
x"00",	-- Hex Addr	410B	16651
x"00",	-- Hex Addr	410C	16652
x"00",	-- Hex Addr	410D	16653
x"00",	-- Hex Addr	410E	16654
x"00",	-- Hex Addr	410F	16655
x"00",	-- Hex Addr	4110	16656
x"00",	-- Hex Addr	4111	16657
x"00",	-- Hex Addr	4112	16658
x"00",	-- Hex Addr	4113	16659
x"00",	-- Hex Addr	4114	16660
x"00",	-- Hex Addr	4115	16661
x"00",	-- Hex Addr	4116	16662
x"00",	-- Hex Addr	4117	16663
x"00",	-- Hex Addr	4118	16664
x"00",	-- Hex Addr	4119	16665
x"00",	-- Hex Addr	411A	16666
x"00",	-- Hex Addr	411B	16667
x"00",	-- Hex Addr	411C	16668
x"00",	-- Hex Addr	411D	16669
x"00",	-- Hex Addr	411E	16670
x"00",	-- Hex Addr	411F	16671
x"00",	-- Hex Addr	4120	16672
x"00",	-- Hex Addr	4121	16673
x"00",	-- Hex Addr	4122	16674
x"00",	-- Hex Addr	4123	16675
x"00",	-- Hex Addr	4124	16676
x"00",	-- Hex Addr	4125	16677
x"00",	-- Hex Addr	4126	16678
x"00",	-- Hex Addr	4127	16679
x"00",	-- Hex Addr	4128	16680
x"00",	-- Hex Addr	4129	16681
x"00",	-- Hex Addr	412A	16682
x"00",	-- Hex Addr	412B	16683
x"00",	-- Hex Addr	412C	16684
x"00",	-- Hex Addr	412D	16685
x"00",	-- Hex Addr	412E	16686
x"00",	-- Hex Addr	412F	16687
x"00",	-- Hex Addr	4130	16688
x"00",	-- Hex Addr	4131	16689
x"00",	-- Hex Addr	4132	16690
x"00",	-- Hex Addr	4133	16691
x"00",	-- Hex Addr	4134	16692
x"00",	-- Hex Addr	4135	16693
x"00",	-- Hex Addr	4136	16694
x"00",	-- Hex Addr	4137	16695
x"00",	-- Hex Addr	4138	16696
x"00",	-- Hex Addr	4139	16697
x"00",	-- Hex Addr	413A	16698
x"00",	-- Hex Addr	413B	16699
x"00",	-- Hex Addr	413C	16700
x"00",	-- Hex Addr	413D	16701
x"00",	-- Hex Addr	413E	16702
x"00",	-- Hex Addr	413F	16703
x"00",	-- Hex Addr	4140	16704
x"00",	-- Hex Addr	4141	16705
x"00",	-- Hex Addr	4142	16706
x"00",	-- Hex Addr	4143	16707
x"00",	-- Hex Addr	4144	16708
x"00",	-- Hex Addr	4145	16709
x"00",	-- Hex Addr	4146	16710
x"00",	-- Hex Addr	4147	16711
x"00",	-- Hex Addr	4148	16712
x"00",	-- Hex Addr	4149	16713
x"00",	-- Hex Addr	414A	16714
x"00",	-- Hex Addr	414B	16715
x"00",	-- Hex Addr	414C	16716
x"00",	-- Hex Addr	414D	16717
x"00",	-- Hex Addr	414E	16718
x"00",	-- Hex Addr	414F	16719
x"00",	-- Hex Addr	4150	16720
x"00",	-- Hex Addr	4151	16721
x"00",	-- Hex Addr	4152	16722
x"00",	-- Hex Addr	4153	16723
x"00",	-- Hex Addr	4154	16724
x"00",	-- Hex Addr	4155	16725
x"00",	-- Hex Addr	4156	16726
x"00",	-- Hex Addr	4157	16727
x"00",	-- Hex Addr	4158	16728
x"00",	-- Hex Addr	4159	16729
x"00",	-- Hex Addr	415A	16730
x"00",	-- Hex Addr	415B	16731
x"00",	-- Hex Addr	415C	16732
x"00",	-- Hex Addr	415D	16733
x"00",	-- Hex Addr	415E	16734
x"00",	-- Hex Addr	415F	16735
x"00",	-- Hex Addr	4160	16736
x"00",	-- Hex Addr	4161	16737
x"00",	-- Hex Addr	4162	16738
x"00",	-- Hex Addr	4163	16739
x"00",	-- Hex Addr	4164	16740
x"00",	-- Hex Addr	4165	16741
x"00",	-- Hex Addr	4166	16742
x"00",	-- Hex Addr	4167	16743
x"00",	-- Hex Addr	4168	16744
x"00",	-- Hex Addr	4169	16745
x"00",	-- Hex Addr	416A	16746
x"00",	-- Hex Addr	416B	16747
x"00",	-- Hex Addr	416C	16748
x"00",	-- Hex Addr	416D	16749
x"00",	-- Hex Addr	416E	16750
x"00",	-- Hex Addr	416F	16751
x"00",	-- Hex Addr	4170	16752
x"00",	-- Hex Addr	4171	16753
x"00",	-- Hex Addr	4172	16754
x"00",	-- Hex Addr	4173	16755
x"00",	-- Hex Addr	4174	16756
x"00",	-- Hex Addr	4175	16757
x"00",	-- Hex Addr	4176	16758
x"00",	-- Hex Addr	4177	16759
x"00",	-- Hex Addr	4178	16760
x"00",	-- Hex Addr	4179	16761
x"00",	-- Hex Addr	417A	16762
x"00",	-- Hex Addr	417B	16763
x"00",	-- Hex Addr	417C	16764
x"00",	-- Hex Addr	417D	16765
x"00",	-- Hex Addr	417E	16766
x"00",	-- Hex Addr	417F	16767
x"00",	-- Hex Addr	4180	16768
x"00",	-- Hex Addr	4181	16769
x"00",	-- Hex Addr	4182	16770
x"00",	-- Hex Addr	4183	16771
x"00",	-- Hex Addr	4184	16772
x"00",	-- Hex Addr	4185	16773
x"00",	-- Hex Addr	4186	16774
x"00",	-- Hex Addr	4187	16775
x"00",	-- Hex Addr	4188	16776
x"00",	-- Hex Addr	4189	16777
x"00",	-- Hex Addr	418A	16778
x"00",	-- Hex Addr	418B	16779
x"00",	-- Hex Addr	418C	16780
x"00",	-- Hex Addr	418D	16781
x"00",	-- Hex Addr	418E	16782
x"00",	-- Hex Addr	418F	16783
x"00",	-- Hex Addr	4190	16784
x"00",	-- Hex Addr	4191	16785
x"00",	-- Hex Addr	4192	16786
x"00",	-- Hex Addr	4193	16787
x"00",	-- Hex Addr	4194	16788
x"00",	-- Hex Addr	4195	16789
x"00",	-- Hex Addr	4196	16790
x"00",	-- Hex Addr	4197	16791
x"00",	-- Hex Addr	4198	16792
x"00",	-- Hex Addr	4199	16793
x"00",	-- Hex Addr	419A	16794
x"00",	-- Hex Addr	419B	16795
x"00",	-- Hex Addr	419C	16796
x"00",	-- Hex Addr	419D	16797
x"00",	-- Hex Addr	419E	16798
x"00",	-- Hex Addr	419F	16799
x"00",	-- Hex Addr	41A0	16800
x"00",	-- Hex Addr	41A1	16801
x"00",	-- Hex Addr	41A2	16802
x"00",	-- Hex Addr	41A3	16803
x"00",	-- Hex Addr	41A4	16804
x"00",	-- Hex Addr	41A5	16805
x"00",	-- Hex Addr	41A6	16806
x"00",	-- Hex Addr	41A7	16807
x"00",	-- Hex Addr	41A8	16808
x"00",	-- Hex Addr	41A9	16809
x"00",	-- Hex Addr	41AA	16810
x"00",	-- Hex Addr	41AB	16811
x"00",	-- Hex Addr	41AC	16812
x"00",	-- Hex Addr	41AD	16813
x"00",	-- Hex Addr	41AE	16814
x"00",	-- Hex Addr	41AF	16815
x"00",	-- Hex Addr	41B0	16816
x"00",	-- Hex Addr	41B1	16817
x"00",	-- Hex Addr	41B2	16818
x"00",	-- Hex Addr	41B3	16819
x"00",	-- Hex Addr	41B4	16820
x"00",	-- Hex Addr	41B5	16821
x"00",	-- Hex Addr	41B6	16822
x"00",	-- Hex Addr	41B7	16823
x"00",	-- Hex Addr	41B8	16824
x"00",	-- Hex Addr	41B9	16825
x"00",	-- Hex Addr	41BA	16826
x"00",	-- Hex Addr	41BB	16827
x"00",	-- Hex Addr	41BC	16828
x"00",	-- Hex Addr	41BD	16829
x"00",	-- Hex Addr	41BE	16830
x"00",	-- Hex Addr	41BF	16831
x"00",	-- Hex Addr	41C0	16832
x"00",	-- Hex Addr	41C1	16833
x"00",	-- Hex Addr	41C2	16834
x"00",	-- Hex Addr	41C3	16835
x"00",	-- Hex Addr	41C4	16836
x"00",	-- Hex Addr	41C5	16837
x"00",	-- Hex Addr	41C6	16838
x"00",	-- Hex Addr	41C7	16839
x"00",	-- Hex Addr	41C8	16840
x"00",	-- Hex Addr	41C9	16841
x"00",	-- Hex Addr	41CA	16842
x"00",	-- Hex Addr	41CB	16843
x"00",	-- Hex Addr	41CC	16844
x"00",	-- Hex Addr	41CD	16845
x"00",	-- Hex Addr	41CE	16846
x"00",	-- Hex Addr	41CF	16847
x"00",	-- Hex Addr	41D0	16848
x"00",	-- Hex Addr	41D1	16849
x"00",	-- Hex Addr	41D2	16850
x"00",	-- Hex Addr	41D3	16851
x"00",	-- Hex Addr	41D4	16852
x"00",	-- Hex Addr	41D5	16853
x"00",	-- Hex Addr	41D6	16854
x"00",	-- Hex Addr	41D7	16855
x"00",	-- Hex Addr	41D8	16856
x"00",	-- Hex Addr	41D9	16857
x"00",	-- Hex Addr	41DA	16858
x"00",	-- Hex Addr	41DB	16859
x"00",	-- Hex Addr	41DC	16860
x"00",	-- Hex Addr	41DD	16861
x"00",	-- Hex Addr	41DE	16862
x"00",	-- Hex Addr	41DF	16863
x"00",	-- Hex Addr	41E0	16864
x"00",	-- Hex Addr	41E1	16865
x"00",	-- Hex Addr	41E2	16866
x"00",	-- Hex Addr	41E3	16867
x"00",	-- Hex Addr	41E4	16868
x"00",	-- Hex Addr	41E5	16869
x"00",	-- Hex Addr	41E6	16870
x"00",	-- Hex Addr	41E7	16871
x"00",	-- Hex Addr	41E8	16872
x"00",	-- Hex Addr	41E9	16873
x"00",	-- Hex Addr	41EA	16874
x"00",	-- Hex Addr	41EB	16875
x"00",	-- Hex Addr	41EC	16876
x"00",	-- Hex Addr	41ED	16877
x"00",	-- Hex Addr	41EE	16878
x"00",	-- Hex Addr	41EF	16879
x"00",	-- Hex Addr	41F0	16880
x"00",	-- Hex Addr	41F1	16881
x"00",	-- Hex Addr	41F2	16882
x"00",	-- Hex Addr	41F3	16883
x"00",	-- Hex Addr	41F4	16884
x"00",	-- Hex Addr	41F5	16885
x"00",	-- Hex Addr	41F6	16886
x"00",	-- Hex Addr	41F7	16887
x"00",	-- Hex Addr	41F8	16888
x"00",	-- Hex Addr	41F9	16889
x"00",	-- Hex Addr	41FA	16890
x"00",	-- Hex Addr	41FB	16891
x"00",	-- Hex Addr	41FC	16892
x"00",	-- Hex Addr	41FD	16893
x"00",	-- Hex Addr	41FE	16894
x"00",	-- Hex Addr	41FF	16895
x"00",	-- Hex Addr	4200	16896
x"00",	-- Hex Addr	4201	16897
x"00",	-- Hex Addr	4202	16898
x"00",	-- Hex Addr	4203	16899
x"00",	-- Hex Addr	4204	16900
x"00",	-- Hex Addr	4205	16901
x"00",	-- Hex Addr	4206	16902
x"00",	-- Hex Addr	4207	16903
x"00",	-- Hex Addr	4208	16904
x"00",	-- Hex Addr	4209	16905
x"00",	-- Hex Addr	420A	16906
x"00",	-- Hex Addr	420B	16907
x"00",	-- Hex Addr	420C	16908
x"00",	-- Hex Addr	420D	16909
x"00",	-- Hex Addr	420E	16910
x"00",	-- Hex Addr	420F	16911
x"00",	-- Hex Addr	4210	16912
x"00",	-- Hex Addr	4211	16913
x"00",	-- Hex Addr	4212	16914
x"00",	-- Hex Addr	4213	16915
x"00",	-- Hex Addr	4214	16916
x"00",	-- Hex Addr	4215	16917
x"00",	-- Hex Addr	4216	16918
x"00",	-- Hex Addr	4217	16919
x"00",	-- Hex Addr	4218	16920
x"00",	-- Hex Addr	4219	16921
x"00",	-- Hex Addr	421A	16922
x"00",	-- Hex Addr	421B	16923
x"00",	-- Hex Addr	421C	16924
x"00",	-- Hex Addr	421D	16925
x"00",	-- Hex Addr	421E	16926
x"00",	-- Hex Addr	421F	16927
x"00",	-- Hex Addr	4220	16928
x"00",	-- Hex Addr	4221	16929
x"00",	-- Hex Addr	4222	16930
x"00",	-- Hex Addr	4223	16931
x"00",	-- Hex Addr	4224	16932
x"00",	-- Hex Addr	4225	16933
x"00",	-- Hex Addr	4226	16934
x"00",	-- Hex Addr	4227	16935
x"00",	-- Hex Addr	4228	16936
x"00",	-- Hex Addr	4229	16937
x"00",	-- Hex Addr	422A	16938
x"00",	-- Hex Addr	422B	16939
x"00",	-- Hex Addr	422C	16940
x"00",	-- Hex Addr	422D	16941
x"00",	-- Hex Addr	422E	16942
x"00",	-- Hex Addr	422F	16943
x"00",	-- Hex Addr	4230	16944
x"00",	-- Hex Addr	4231	16945
x"00",	-- Hex Addr	4232	16946
x"00",	-- Hex Addr	4233	16947
x"00",	-- Hex Addr	4234	16948
x"00",	-- Hex Addr	4235	16949
x"00",	-- Hex Addr	4236	16950
x"00",	-- Hex Addr	4237	16951
x"00",	-- Hex Addr	4238	16952
x"00",	-- Hex Addr	4239	16953
x"00",	-- Hex Addr	423A	16954
x"00",	-- Hex Addr	423B	16955
x"00",	-- Hex Addr	423C	16956
x"00",	-- Hex Addr	423D	16957
x"00",	-- Hex Addr	423E	16958
x"00",	-- Hex Addr	423F	16959
x"00",	-- Hex Addr	4240	16960
x"00",	-- Hex Addr	4241	16961
x"00",	-- Hex Addr	4242	16962
x"00",	-- Hex Addr	4243	16963
x"00",	-- Hex Addr	4244	16964
x"00",	-- Hex Addr	4245	16965
x"00",	-- Hex Addr	4246	16966
x"00",	-- Hex Addr	4247	16967
x"00",	-- Hex Addr	4248	16968
x"00",	-- Hex Addr	4249	16969
x"00",	-- Hex Addr	424A	16970
x"00",	-- Hex Addr	424B	16971
x"00",	-- Hex Addr	424C	16972
x"00",	-- Hex Addr	424D	16973
x"00",	-- Hex Addr	424E	16974
x"00",	-- Hex Addr	424F	16975
x"00",	-- Hex Addr	4250	16976
x"00",	-- Hex Addr	4251	16977
x"00",	-- Hex Addr	4252	16978
x"00",	-- Hex Addr	4253	16979
x"00",	-- Hex Addr	4254	16980
x"00",	-- Hex Addr	4255	16981
x"00",	-- Hex Addr	4256	16982
x"00",	-- Hex Addr	4257	16983
x"00",	-- Hex Addr	4258	16984
x"00",	-- Hex Addr	4259	16985
x"00",	-- Hex Addr	425A	16986
x"00",	-- Hex Addr	425B	16987
x"00",	-- Hex Addr	425C	16988
x"00",	-- Hex Addr	425D	16989
x"00",	-- Hex Addr	425E	16990
x"00",	-- Hex Addr	425F	16991
x"00",	-- Hex Addr	4260	16992
x"00",	-- Hex Addr	4261	16993
x"00",	-- Hex Addr	4262	16994
x"00",	-- Hex Addr	4263	16995
x"00",	-- Hex Addr	4264	16996
x"00",	-- Hex Addr	4265	16997
x"00",	-- Hex Addr	4266	16998
x"00",	-- Hex Addr	4267	16999
x"00",	-- Hex Addr	4268	17000
x"00",	-- Hex Addr	4269	17001
x"00",	-- Hex Addr	426A	17002
x"00",	-- Hex Addr	426B	17003
x"00",	-- Hex Addr	426C	17004
x"00",	-- Hex Addr	426D	17005
x"00",	-- Hex Addr	426E	17006
x"00",	-- Hex Addr	426F	17007
x"00",	-- Hex Addr	4270	17008
x"00",	-- Hex Addr	4271	17009
x"00",	-- Hex Addr	4272	17010
x"00",	-- Hex Addr	4273	17011
x"00",	-- Hex Addr	4274	17012
x"00",	-- Hex Addr	4275	17013
x"00",	-- Hex Addr	4276	17014
x"00",	-- Hex Addr	4277	17015
x"00",	-- Hex Addr	4278	17016
x"00",	-- Hex Addr	4279	17017
x"00",	-- Hex Addr	427A	17018
x"00",	-- Hex Addr	427B	17019
x"00",	-- Hex Addr	427C	17020
x"00",	-- Hex Addr	427D	17021
x"00",	-- Hex Addr	427E	17022
x"00",	-- Hex Addr	427F	17023
x"00",	-- Hex Addr	4280	17024
x"00",	-- Hex Addr	4281	17025
x"00",	-- Hex Addr	4282	17026
x"00",	-- Hex Addr	4283	17027
x"00",	-- Hex Addr	4284	17028
x"00",	-- Hex Addr	4285	17029
x"00",	-- Hex Addr	4286	17030
x"00",	-- Hex Addr	4287	17031
x"00",	-- Hex Addr	4288	17032
x"00",	-- Hex Addr	4289	17033
x"00",	-- Hex Addr	428A	17034
x"00",	-- Hex Addr	428B	17035
x"00",	-- Hex Addr	428C	17036
x"00",	-- Hex Addr	428D	17037
x"00",	-- Hex Addr	428E	17038
x"00",	-- Hex Addr	428F	17039
x"00",	-- Hex Addr	4290	17040
x"00",	-- Hex Addr	4291	17041
x"00",	-- Hex Addr	4292	17042
x"00",	-- Hex Addr	4293	17043
x"00",	-- Hex Addr	4294	17044
x"00",	-- Hex Addr	4295	17045
x"00",	-- Hex Addr	4296	17046
x"00",	-- Hex Addr	4297	17047
x"00",	-- Hex Addr	4298	17048
x"00",	-- Hex Addr	4299	17049
x"00",	-- Hex Addr	429A	17050
x"00",	-- Hex Addr	429B	17051
x"00",	-- Hex Addr	429C	17052
x"00",	-- Hex Addr	429D	17053
x"00",	-- Hex Addr	429E	17054
x"00",	-- Hex Addr	429F	17055
x"00",	-- Hex Addr	42A0	17056
x"00",	-- Hex Addr	42A1	17057
x"00",	-- Hex Addr	42A2	17058
x"00",	-- Hex Addr	42A3	17059
x"00",	-- Hex Addr	42A4	17060
x"00",	-- Hex Addr	42A5	17061
x"00",	-- Hex Addr	42A6	17062
x"00",	-- Hex Addr	42A7	17063
x"00",	-- Hex Addr	42A8	17064
x"00",	-- Hex Addr	42A9	17065
x"00",	-- Hex Addr	42AA	17066
x"00",	-- Hex Addr	42AB	17067
x"00",	-- Hex Addr	42AC	17068
x"00",	-- Hex Addr	42AD	17069
x"00",	-- Hex Addr	42AE	17070
x"00",	-- Hex Addr	42AF	17071
x"00",	-- Hex Addr	42B0	17072
x"00",	-- Hex Addr	42B1	17073
x"00",	-- Hex Addr	42B2	17074
x"00",	-- Hex Addr	42B3	17075
x"00",	-- Hex Addr	42B4	17076
x"00",	-- Hex Addr	42B5	17077
x"00",	-- Hex Addr	42B6	17078
x"00",	-- Hex Addr	42B7	17079
x"00",	-- Hex Addr	42B8	17080
x"00",	-- Hex Addr	42B9	17081
x"00",	-- Hex Addr	42BA	17082
x"00",	-- Hex Addr	42BB	17083
x"00",	-- Hex Addr	42BC	17084
x"00",	-- Hex Addr	42BD	17085
x"00",	-- Hex Addr	42BE	17086
x"00",	-- Hex Addr	42BF	17087
x"00",	-- Hex Addr	42C0	17088
x"00",	-- Hex Addr	42C1	17089
x"00",	-- Hex Addr	42C2	17090
x"00",	-- Hex Addr	42C3	17091
x"00",	-- Hex Addr	42C4	17092
x"00",	-- Hex Addr	42C5	17093
x"00",	-- Hex Addr	42C6	17094
x"00",	-- Hex Addr	42C7	17095
x"00",	-- Hex Addr	42C8	17096
x"00",	-- Hex Addr	42C9	17097
x"00",	-- Hex Addr	42CA	17098
x"00",	-- Hex Addr	42CB	17099
x"00",	-- Hex Addr	42CC	17100
x"00",	-- Hex Addr	42CD	17101
x"00",	-- Hex Addr	42CE	17102
x"00",	-- Hex Addr	42CF	17103
x"00",	-- Hex Addr	42D0	17104
x"00",	-- Hex Addr	42D1	17105
x"00",	-- Hex Addr	42D2	17106
x"00",	-- Hex Addr	42D3	17107
x"00",	-- Hex Addr	42D4	17108
x"00",	-- Hex Addr	42D5	17109
x"00",	-- Hex Addr	42D6	17110
x"00",	-- Hex Addr	42D7	17111
x"00",	-- Hex Addr	42D8	17112
x"00",	-- Hex Addr	42D9	17113
x"00",	-- Hex Addr	42DA	17114
x"00",	-- Hex Addr	42DB	17115
x"00",	-- Hex Addr	42DC	17116
x"00",	-- Hex Addr	42DD	17117
x"00",	-- Hex Addr	42DE	17118
x"00",	-- Hex Addr	42DF	17119
x"00",	-- Hex Addr	42E0	17120
x"00",	-- Hex Addr	42E1	17121
x"00",	-- Hex Addr	42E2	17122
x"00",	-- Hex Addr	42E3	17123
x"00",	-- Hex Addr	42E4	17124
x"00",	-- Hex Addr	42E5	17125
x"00",	-- Hex Addr	42E6	17126
x"00",	-- Hex Addr	42E7	17127
x"00",	-- Hex Addr	42E8	17128
x"00",	-- Hex Addr	42E9	17129
x"00",	-- Hex Addr	42EA	17130
x"00",	-- Hex Addr	42EB	17131
x"00",	-- Hex Addr	42EC	17132
x"00",	-- Hex Addr	42ED	17133
x"00",	-- Hex Addr	42EE	17134
x"00",	-- Hex Addr	42EF	17135
x"00",	-- Hex Addr	42F0	17136
x"00",	-- Hex Addr	42F1	17137
x"00",	-- Hex Addr	42F2	17138
x"00",	-- Hex Addr	42F3	17139
x"00",	-- Hex Addr	42F4	17140
x"00",	-- Hex Addr	42F5	17141
x"00",	-- Hex Addr	42F6	17142
x"00",	-- Hex Addr	42F7	17143
x"00",	-- Hex Addr	42F8	17144
x"00",	-- Hex Addr	42F9	17145
x"00",	-- Hex Addr	42FA	17146
x"00",	-- Hex Addr	42FB	17147
x"00",	-- Hex Addr	42FC	17148
x"00",	-- Hex Addr	42FD	17149
x"00",	-- Hex Addr	42FE	17150
x"00",	-- Hex Addr	42FF	17151
x"00",	-- Hex Addr	4300	17152
x"00",	-- Hex Addr	4301	17153
x"00",	-- Hex Addr	4302	17154
x"00",	-- Hex Addr	4303	17155
x"00",	-- Hex Addr	4304	17156
x"00",	-- Hex Addr	4305	17157
x"00",	-- Hex Addr	4306	17158
x"00",	-- Hex Addr	4307	17159
x"00",	-- Hex Addr	4308	17160
x"00",	-- Hex Addr	4309	17161
x"00",	-- Hex Addr	430A	17162
x"00",	-- Hex Addr	430B	17163
x"00",	-- Hex Addr	430C	17164
x"00",	-- Hex Addr	430D	17165
x"00",	-- Hex Addr	430E	17166
x"00",	-- Hex Addr	430F	17167
x"00",	-- Hex Addr	4310	17168
x"00",	-- Hex Addr	4311	17169
x"00",	-- Hex Addr	4312	17170
x"00",	-- Hex Addr	4313	17171
x"00",	-- Hex Addr	4314	17172
x"00",	-- Hex Addr	4315	17173
x"00",	-- Hex Addr	4316	17174
x"00",	-- Hex Addr	4317	17175
x"00",	-- Hex Addr	4318	17176
x"00",	-- Hex Addr	4319	17177
x"00",	-- Hex Addr	431A	17178
x"00",	-- Hex Addr	431B	17179
x"00",	-- Hex Addr	431C	17180
x"00",	-- Hex Addr	431D	17181
x"00",	-- Hex Addr	431E	17182
x"00",	-- Hex Addr	431F	17183
x"00",	-- Hex Addr	4320	17184
x"00",	-- Hex Addr	4321	17185
x"00",	-- Hex Addr	4322	17186
x"00",	-- Hex Addr	4323	17187
x"00",	-- Hex Addr	4324	17188
x"00",	-- Hex Addr	4325	17189
x"00",	-- Hex Addr	4326	17190
x"00",	-- Hex Addr	4327	17191
x"00",	-- Hex Addr	4328	17192
x"00",	-- Hex Addr	4329	17193
x"00",	-- Hex Addr	432A	17194
x"00",	-- Hex Addr	432B	17195
x"00",	-- Hex Addr	432C	17196
x"00",	-- Hex Addr	432D	17197
x"00",	-- Hex Addr	432E	17198
x"00",	-- Hex Addr	432F	17199
x"00",	-- Hex Addr	4330	17200
x"00",	-- Hex Addr	4331	17201
x"00",	-- Hex Addr	4332	17202
x"00",	-- Hex Addr	4333	17203
x"00",	-- Hex Addr	4334	17204
x"00",	-- Hex Addr	4335	17205
x"00",	-- Hex Addr	4336	17206
x"00",	-- Hex Addr	4337	17207
x"00",	-- Hex Addr	4338	17208
x"00",	-- Hex Addr	4339	17209
x"00",	-- Hex Addr	433A	17210
x"00",	-- Hex Addr	433B	17211
x"00",	-- Hex Addr	433C	17212
x"00",	-- Hex Addr	433D	17213
x"00",	-- Hex Addr	433E	17214
x"00",	-- Hex Addr	433F	17215
x"00",	-- Hex Addr	4340	17216
x"00",	-- Hex Addr	4341	17217
x"00",	-- Hex Addr	4342	17218
x"00",	-- Hex Addr	4343	17219
x"00",	-- Hex Addr	4344	17220
x"00",	-- Hex Addr	4345	17221
x"00",	-- Hex Addr	4346	17222
x"00",	-- Hex Addr	4347	17223
x"00",	-- Hex Addr	4348	17224
x"00",	-- Hex Addr	4349	17225
x"00",	-- Hex Addr	434A	17226
x"00",	-- Hex Addr	434B	17227
x"00",	-- Hex Addr	434C	17228
x"00",	-- Hex Addr	434D	17229
x"00",	-- Hex Addr	434E	17230
x"00",	-- Hex Addr	434F	17231
x"00",	-- Hex Addr	4350	17232
x"00",	-- Hex Addr	4351	17233
x"00",	-- Hex Addr	4352	17234
x"00",	-- Hex Addr	4353	17235
x"00",	-- Hex Addr	4354	17236
x"00",	-- Hex Addr	4355	17237
x"00",	-- Hex Addr	4356	17238
x"00",	-- Hex Addr	4357	17239
x"00",	-- Hex Addr	4358	17240
x"00",	-- Hex Addr	4359	17241
x"00",	-- Hex Addr	435A	17242
x"00",	-- Hex Addr	435B	17243
x"00",	-- Hex Addr	435C	17244
x"00",	-- Hex Addr	435D	17245
x"00",	-- Hex Addr	435E	17246
x"00",	-- Hex Addr	435F	17247
x"00",	-- Hex Addr	4360	17248
x"00",	-- Hex Addr	4361	17249
x"00",	-- Hex Addr	4362	17250
x"00",	-- Hex Addr	4363	17251
x"00",	-- Hex Addr	4364	17252
x"00",	-- Hex Addr	4365	17253
x"00",	-- Hex Addr	4366	17254
x"00",	-- Hex Addr	4367	17255
x"00",	-- Hex Addr	4368	17256
x"00",	-- Hex Addr	4369	17257
x"00",	-- Hex Addr	436A	17258
x"00",	-- Hex Addr	436B	17259
x"00",	-- Hex Addr	436C	17260
x"00",	-- Hex Addr	436D	17261
x"00",	-- Hex Addr	436E	17262
x"00",	-- Hex Addr	436F	17263
x"00",	-- Hex Addr	4370	17264
x"00",	-- Hex Addr	4371	17265
x"00",	-- Hex Addr	4372	17266
x"00",	-- Hex Addr	4373	17267
x"00",	-- Hex Addr	4374	17268
x"00",	-- Hex Addr	4375	17269
x"00",	-- Hex Addr	4376	17270
x"00",	-- Hex Addr	4377	17271
x"00",	-- Hex Addr	4378	17272
x"00",	-- Hex Addr	4379	17273
x"00",	-- Hex Addr	437A	17274
x"00",	-- Hex Addr	437B	17275
x"00",	-- Hex Addr	437C	17276
x"00",	-- Hex Addr	437D	17277
x"00",	-- Hex Addr	437E	17278
x"00",	-- Hex Addr	437F	17279
x"00",	-- Hex Addr	4380	17280
x"00",	-- Hex Addr	4381	17281
x"00",	-- Hex Addr	4382	17282
x"00",	-- Hex Addr	4383	17283
x"00",	-- Hex Addr	4384	17284
x"00",	-- Hex Addr	4385	17285
x"00",	-- Hex Addr	4386	17286
x"00",	-- Hex Addr	4387	17287
x"00",	-- Hex Addr	4388	17288
x"00",	-- Hex Addr	4389	17289
x"00",	-- Hex Addr	438A	17290
x"00",	-- Hex Addr	438B	17291
x"00",	-- Hex Addr	438C	17292
x"00",	-- Hex Addr	438D	17293
x"00",	-- Hex Addr	438E	17294
x"00",	-- Hex Addr	438F	17295
x"00",	-- Hex Addr	4390	17296
x"00",	-- Hex Addr	4391	17297
x"00",	-- Hex Addr	4392	17298
x"00",	-- Hex Addr	4393	17299
x"00",	-- Hex Addr	4394	17300
x"00",	-- Hex Addr	4395	17301
x"00",	-- Hex Addr	4396	17302
x"00",	-- Hex Addr	4397	17303
x"00",	-- Hex Addr	4398	17304
x"00",	-- Hex Addr	4399	17305
x"00",	-- Hex Addr	439A	17306
x"00",	-- Hex Addr	439B	17307
x"00",	-- Hex Addr	439C	17308
x"00",	-- Hex Addr	439D	17309
x"00",	-- Hex Addr	439E	17310
x"00",	-- Hex Addr	439F	17311
x"00",	-- Hex Addr	43A0	17312
x"00",	-- Hex Addr	43A1	17313
x"00",	-- Hex Addr	43A2	17314
x"00",	-- Hex Addr	43A3	17315
x"00",	-- Hex Addr	43A4	17316
x"00",	-- Hex Addr	43A5	17317
x"00",	-- Hex Addr	43A6	17318
x"00",	-- Hex Addr	43A7	17319
x"00",	-- Hex Addr	43A8	17320
x"00",	-- Hex Addr	43A9	17321
x"00",	-- Hex Addr	43AA	17322
x"00",	-- Hex Addr	43AB	17323
x"00",	-- Hex Addr	43AC	17324
x"00",	-- Hex Addr	43AD	17325
x"00",	-- Hex Addr	43AE	17326
x"00",	-- Hex Addr	43AF	17327
x"00",	-- Hex Addr	43B0	17328
x"00",	-- Hex Addr	43B1	17329
x"00",	-- Hex Addr	43B2	17330
x"00",	-- Hex Addr	43B3	17331
x"00",	-- Hex Addr	43B4	17332
x"00",	-- Hex Addr	43B5	17333
x"00",	-- Hex Addr	43B6	17334
x"00",	-- Hex Addr	43B7	17335
x"00",	-- Hex Addr	43B8	17336
x"00",	-- Hex Addr	43B9	17337
x"00",	-- Hex Addr	43BA	17338
x"00",	-- Hex Addr	43BB	17339
x"00",	-- Hex Addr	43BC	17340
x"00",	-- Hex Addr	43BD	17341
x"00",	-- Hex Addr	43BE	17342
x"00",	-- Hex Addr	43BF	17343
x"00",	-- Hex Addr	43C0	17344
x"00",	-- Hex Addr	43C1	17345
x"00",	-- Hex Addr	43C2	17346
x"00",	-- Hex Addr	43C3	17347
x"00",	-- Hex Addr	43C4	17348
x"00",	-- Hex Addr	43C5	17349
x"00",	-- Hex Addr	43C6	17350
x"00",	-- Hex Addr	43C7	17351
x"00",	-- Hex Addr	43C8	17352
x"00",	-- Hex Addr	43C9	17353
x"00",	-- Hex Addr	43CA	17354
x"00",	-- Hex Addr	43CB	17355
x"00",	-- Hex Addr	43CC	17356
x"00",	-- Hex Addr	43CD	17357
x"00",	-- Hex Addr	43CE	17358
x"00",	-- Hex Addr	43CF	17359
x"00",	-- Hex Addr	43D0	17360
x"00",	-- Hex Addr	43D1	17361
x"00",	-- Hex Addr	43D2	17362
x"00",	-- Hex Addr	43D3	17363
x"00",	-- Hex Addr	43D4	17364
x"00",	-- Hex Addr	43D5	17365
x"00",	-- Hex Addr	43D6	17366
x"00",	-- Hex Addr	43D7	17367
x"00",	-- Hex Addr	43D8	17368
x"00",	-- Hex Addr	43D9	17369
x"00",	-- Hex Addr	43DA	17370
x"00",	-- Hex Addr	43DB	17371
x"00",	-- Hex Addr	43DC	17372
x"00",	-- Hex Addr	43DD	17373
x"00",	-- Hex Addr	43DE	17374
x"00",	-- Hex Addr	43DF	17375
x"00",	-- Hex Addr	43E0	17376
x"00",	-- Hex Addr	43E1	17377
x"00",	-- Hex Addr	43E2	17378
x"00",	-- Hex Addr	43E3	17379
x"00",	-- Hex Addr	43E4	17380
x"00",	-- Hex Addr	43E5	17381
x"00",	-- Hex Addr	43E6	17382
x"00",	-- Hex Addr	43E7	17383
x"00",	-- Hex Addr	43E8	17384
x"00",	-- Hex Addr	43E9	17385
x"00",	-- Hex Addr	43EA	17386
x"00",	-- Hex Addr	43EB	17387
x"00",	-- Hex Addr	43EC	17388
x"00",	-- Hex Addr	43ED	17389
x"00",	-- Hex Addr	43EE	17390
x"00",	-- Hex Addr	43EF	17391
x"00",	-- Hex Addr	43F0	17392
x"00",	-- Hex Addr	43F1	17393
x"00",	-- Hex Addr	43F2	17394
x"00",	-- Hex Addr	43F3	17395
x"00",	-- Hex Addr	43F4	17396
x"00",	-- Hex Addr	43F5	17397
x"00",	-- Hex Addr	43F6	17398
x"00",	-- Hex Addr	43F7	17399
x"00",	-- Hex Addr	43F8	17400
x"00",	-- Hex Addr	43F9	17401
x"00",	-- Hex Addr	43FA	17402
x"00",	-- Hex Addr	43FB	17403
x"00",	-- Hex Addr	43FC	17404
x"00",	-- Hex Addr	43FD	17405
x"00",	-- Hex Addr	43FE	17406
x"00",	-- Hex Addr	43FF	17407
x"00",	-- Hex Addr	4400	17408
x"00",	-- Hex Addr	4401	17409
x"00",	-- Hex Addr	4402	17410
x"00",	-- Hex Addr	4403	17411
x"00",	-- Hex Addr	4404	17412
x"00",	-- Hex Addr	4405	17413
x"00",	-- Hex Addr	4406	17414
x"00",	-- Hex Addr	4407	17415
x"00",	-- Hex Addr	4408	17416
x"00",	-- Hex Addr	4409	17417
x"00",	-- Hex Addr	440A	17418
x"00",	-- Hex Addr	440B	17419
x"00",	-- Hex Addr	440C	17420
x"00",	-- Hex Addr	440D	17421
x"00",	-- Hex Addr	440E	17422
x"00",	-- Hex Addr	440F	17423
x"00",	-- Hex Addr	4410	17424
x"00",	-- Hex Addr	4411	17425
x"00",	-- Hex Addr	4412	17426
x"00",	-- Hex Addr	4413	17427
x"00",	-- Hex Addr	4414	17428
x"00",	-- Hex Addr	4415	17429
x"00",	-- Hex Addr	4416	17430
x"00",	-- Hex Addr	4417	17431
x"00",	-- Hex Addr	4418	17432
x"00",	-- Hex Addr	4419	17433
x"00",	-- Hex Addr	441A	17434
x"00",	-- Hex Addr	441B	17435
x"00",	-- Hex Addr	441C	17436
x"00",	-- Hex Addr	441D	17437
x"00",	-- Hex Addr	441E	17438
x"00",	-- Hex Addr	441F	17439
x"00",	-- Hex Addr	4420	17440
x"00",	-- Hex Addr	4421	17441
x"00",	-- Hex Addr	4422	17442
x"00",	-- Hex Addr	4423	17443
x"00",	-- Hex Addr	4424	17444
x"00",	-- Hex Addr	4425	17445
x"00",	-- Hex Addr	4426	17446
x"00",	-- Hex Addr	4427	17447
x"00",	-- Hex Addr	4428	17448
x"00",	-- Hex Addr	4429	17449
x"00",	-- Hex Addr	442A	17450
x"00",	-- Hex Addr	442B	17451
x"00",	-- Hex Addr	442C	17452
x"00",	-- Hex Addr	442D	17453
x"00",	-- Hex Addr	442E	17454
x"00",	-- Hex Addr	442F	17455
x"00",	-- Hex Addr	4430	17456
x"00",	-- Hex Addr	4431	17457
x"00",	-- Hex Addr	4432	17458
x"00",	-- Hex Addr	4433	17459
x"00",	-- Hex Addr	4434	17460
x"00",	-- Hex Addr	4435	17461
x"00",	-- Hex Addr	4436	17462
x"00",	-- Hex Addr	4437	17463
x"00",	-- Hex Addr	4438	17464
x"00",	-- Hex Addr	4439	17465
x"00",	-- Hex Addr	443A	17466
x"00",	-- Hex Addr	443B	17467
x"00",	-- Hex Addr	443C	17468
x"00",	-- Hex Addr	443D	17469
x"00",	-- Hex Addr	443E	17470
x"00",	-- Hex Addr	443F	17471
x"00",	-- Hex Addr	4440	17472
x"00",	-- Hex Addr	4441	17473
x"00",	-- Hex Addr	4442	17474
x"00",	-- Hex Addr	4443	17475
x"00",	-- Hex Addr	4444	17476
x"00",	-- Hex Addr	4445	17477
x"00",	-- Hex Addr	4446	17478
x"00",	-- Hex Addr	4447	17479
x"00",	-- Hex Addr	4448	17480
x"00",	-- Hex Addr	4449	17481
x"00",	-- Hex Addr	444A	17482
x"00",	-- Hex Addr	444B	17483
x"00",	-- Hex Addr	444C	17484
x"00",	-- Hex Addr	444D	17485
x"00",	-- Hex Addr	444E	17486
x"00",	-- Hex Addr	444F	17487
x"00",	-- Hex Addr	4450	17488
x"00",	-- Hex Addr	4451	17489
x"00",	-- Hex Addr	4452	17490
x"00",	-- Hex Addr	4453	17491
x"00",	-- Hex Addr	4454	17492
x"00",	-- Hex Addr	4455	17493
x"00",	-- Hex Addr	4456	17494
x"00",	-- Hex Addr	4457	17495
x"00",	-- Hex Addr	4458	17496
x"00",	-- Hex Addr	4459	17497
x"00",	-- Hex Addr	445A	17498
x"00",	-- Hex Addr	445B	17499
x"00",	-- Hex Addr	445C	17500
x"00",	-- Hex Addr	445D	17501
x"00",	-- Hex Addr	445E	17502
x"00",	-- Hex Addr	445F	17503
x"00",	-- Hex Addr	4460	17504
x"00",	-- Hex Addr	4461	17505
x"00",	-- Hex Addr	4462	17506
x"00",	-- Hex Addr	4463	17507
x"00",	-- Hex Addr	4464	17508
x"00",	-- Hex Addr	4465	17509
x"00",	-- Hex Addr	4466	17510
x"00",	-- Hex Addr	4467	17511
x"00",	-- Hex Addr	4468	17512
x"00",	-- Hex Addr	4469	17513
x"00",	-- Hex Addr	446A	17514
x"00",	-- Hex Addr	446B	17515
x"00",	-- Hex Addr	446C	17516
x"00",	-- Hex Addr	446D	17517
x"00",	-- Hex Addr	446E	17518
x"00",	-- Hex Addr	446F	17519
x"00",	-- Hex Addr	4470	17520
x"00",	-- Hex Addr	4471	17521
x"00",	-- Hex Addr	4472	17522
x"00",	-- Hex Addr	4473	17523
x"00",	-- Hex Addr	4474	17524
x"00",	-- Hex Addr	4475	17525
x"00",	-- Hex Addr	4476	17526
x"00",	-- Hex Addr	4477	17527
x"00",	-- Hex Addr	4478	17528
x"00",	-- Hex Addr	4479	17529
x"00",	-- Hex Addr	447A	17530
x"00",	-- Hex Addr	447B	17531
x"00",	-- Hex Addr	447C	17532
x"00",	-- Hex Addr	447D	17533
x"00",	-- Hex Addr	447E	17534
x"00",	-- Hex Addr	447F	17535
x"00",	-- Hex Addr	4480	17536
x"00",	-- Hex Addr	4481	17537
x"00",	-- Hex Addr	4482	17538
x"00",	-- Hex Addr	4483	17539
x"00",	-- Hex Addr	4484	17540
x"00",	-- Hex Addr	4485	17541
x"00",	-- Hex Addr	4486	17542
x"00",	-- Hex Addr	4487	17543
x"00",	-- Hex Addr	4488	17544
x"00",	-- Hex Addr	4489	17545
x"00",	-- Hex Addr	448A	17546
x"00",	-- Hex Addr	448B	17547
x"00",	-- Hex Addr	448C	17548
x"00",	-- Hex Addr	448D	17549
x"00",	-- Hex Addr	448E	17550
x"00",	-- Hex Addr	448F	17551
x"00",	-- Hex Addr	4490	17552
x"00",	-- Hex Addr	4491	17553
x"00",	-- Hex Addr	4492	17554
x"00",	-- Hex Addr	4493	17555
x"00",	-- Hex Addr	4494	17556
x"00",	-- Hex Addr	4495	17557
x"00",	-- Hex Addr	4496	17558
x"00",	-- Hex Addr	4497	17559
x"00",	-- Hex Addr	4498	17560
x"00",	-- Hex Addr	4499	17561
x"00",	-- Hex Addr	449A	17562
x"00",	-- Hex Addr	449B	17563
x"00",	-- Hex Addr	449C	17564
x"00",	-- Hex Addr	449D	17565
x"00",	-- Hex Addr	449E	17566
x"00",	-- Hex Addr	449F	17567
x"00",	-- Hex Addr	44A0	17568
x"00",	-- Hex Addr	44A1	17569
x"00",	-- Hex Addr	44A2	17570
x"00",	-- Hex Addr	44A3	17571
x"00",	-- Hex Addr	44A4	17572
x"00",	-- Hex Addr	44A5	17573
x"00",	-- Hex Addr	44A6	17574
x"00",	-- Hex Addr	44A7	17575
x"00",	-- Hex Addr	44A8	17576
x"00",	-- Hex Addr	44A9	17577
x"00",	-- Hex Addr	44AA	17578
x"00",	-- Hex Addr	44AB	17579
x"00",	-- Hex Addr	44AC	17580
x"00",	-- Hex Addr	44AD	17581
x"00",	-- Hex Addr	44AE	17582
x"00",	-- Hex Addr	44AF	17583
x"00",	-- Hex Addr	44B0	17584
x"00",	-- Hex Addr	44B1	17585
x"00",	-- Hex Addr	44B2	17586
x"00",	-- Hex Addr	44B3	17587
x"00",	-- Hex Addr	44B4	17588
x"00",	-- Hex Addr	44B5	17589
x"00",	-- Hex Addr	44B6	17590
x"00",	-- Hex Addr	44B7	17591
x"00",	-- Hex Addr	44B8	17592
x"00",	-- Hex Addr	44B9	17593
x"00",	-- Hex Addr	44BA	17594
x"00",	-- Hex Addr	44BB	17595
x"00",	-- Hex Addr	44BC	17596
x"00",	-- Hex Addr	44BD	17597
x"00",	-- Hex Addr	44BE	17598
x"00",	-- Hex Addr	44BF	17599
x"00",	-- Hex Addr	44C0	17600
x"00",	-- Hex Addr	44C1	17601
x"00",	-- Hex Addr	44C2	17602
x"00",	-- Hex Addr	44C3	17603
x"00",	-- Hex Addr	44C4	17604
x"00",	-- Hex Addr	44C5	17605
x"00",	-- Hex Addr	44C6	17606
x"00",	-- Hex Addr	44C7	17607
x"00",	-- Hex Addr	44C8	17608
x"00",	-- Hex Addr	44C9	17609
x"00",	-- Hex Addr	44CA	17610
x"00",	-- Hex Addr	44CB	17611
x"00",	-- Hex Addr	44CC	17612
x"00",	-- Hex Addr	44CD	17613
x"00",	-- Hex Addr	44CE	17614
x"00",	-- Hex Addr	44CF	17615
x"00",	-- Hex Addr	44D0	17616
x"00",	-- Hex Addr	44D1	17617
x"00",	-- Hex Addr	44D2	17618
x"00",	-- Hex Addr	44D3	17619
x"00",	-- Hex Addr	44D4	17620
x"00",	-- Hex Addr	44D5	17621
x"00",	-- Hex Addr	44D6	17622
x"00",	-- Hex Addr	44D7	17623
x"00",	-- Hex Addr	44D8	17624
x"00",	-- Hex Addr	44D9	17625
x"00",	-- Hex Addr	44DA	17626
x"00",	-- Hex Addr	44DB	17627
x"00",	-- Hex Addr	44DC	17628
x"00",	-- Hex Addr	44DD	17629
x"00",	-- Hex Addr	44DE	17630
x"00",	-- Hex Addr	44DF	17631
x"00",	-- Hex Addr	44E0	17632
x"00",	-- Hex Addr	44E1	17633
x"00",	-- Hex Addr	44E2	17634
x"00",	-- Hex Addr	44E3	17635
x"00",	-- Hex Addr	44E4	17636
x"00",	-- Hex Addr	44E5	17637
x"00",	-- Hex Addr	44E6	17638
x"00",	-- Hex Addr	44E7	17639
x"00",	-- Hex Addr	44E8	17640
x"00",	-- Hex Addr	44E9	17641
x"00",	-- Hex Addr	44EA	17642
x"00",	-- Hex Addr	44EB	17643
x"00",	-- Hex Addr	44EC	17644
x"00",	-- Hex Addr	44ED	17645
x"00",	-- Hex Addr	44EE	17646
x"00",	-- Hex Addr	44EF	17647
x"00",	-- Hex Addr	44F0	17648
x"00",	-- Hex Addr	44F1	17649
x"00",	-- Hex Addr	44F2	17650
x"00",	-- Hex Addr	44F3	17651
x"00",	-- Hex Addr	44F4	17652
x"00",	-- Hex Addr	44F5	17653
x"00",	-- Hex Addr	44F6	17654
x"00",	-- Hex Addr	44F7	17655
x"00",	-- Hex Addr	44F8	17656
x"00",	-- Hex Addr	44F9	17657
x"00",	-- Hex Addr	44FA	17658
x"00",	-- Hex Addr	44FB	17659
x"00",	-- Hex Addr	44FC	17660
x"00",	-- Hex Addr	44FD	17661
x"00",	-- Hex Addr	44FE	17662
x"00",	-- Hex Addr	44FF	17663
x"00",	-- Hex Addr	4500	17664
x"00",	-- Hex Addr	4501	17665
x"00",	-- Hex Addr	4502	17666
x"00",	-- Hex Addr	4503	17667
x"00",	-- Hex Addr	4504	17668
x"00",	-- Hex Addr	4505	17669
x"00",	-- Hex Addr	4506	17670
x"00",	-- Hex Addr	4507	17671
x"00",	-- Hex Addr	4508	17672
x"00",	-- Hex Addr	4509	17673
x"00",	-- Hex Addr	450A	17674
x"00",	-- Hex Addr	450B	17675
x"00",	-- Hex Addr	450C	17676
x"00",	-- Hex Addr	450D	17677
x"00",	-- Hex Addr	450E	17678
x"00",	-- Hex Addr	450F	17679
x"00",	-- Hex Addr	4510	17680
x"00",	-- Hex Addr	4511	17681
x"00",	-- Hex Addr	4512	17682
x"00",	-- Hex Addr	4513	17683
x"00",	-- Hex Addr	4514	17684
x"00",	-- Hex Addr	4515	17685
x"00",	-- Hex Addr	4516	17686
x"00",	-- Hex Addr	4517	17687
x"00",	-- Hex Addr	4518	17688
x"00",	-- Hex Addr	4519	17689
x"00",	-- Hex Addr	451A	17690
x"00",	-- Hex Addr	451B	17691
x"00",	-- Hex Addr	451C	17692
x"00",	-- Hex Addr	451D	17693
x"00",	-- Hex Addr	451E	17694
x"00",	-- Hex Addr	451F	17695
x"00",	-- Hex Addr	4520	17696
x"00",	-- Hex Addr	4521	17697
x"00",	-- Hex Addr	4522	17698
x"00",	-- Hex Addr	4523	17699
x"00",	-- Hex Addr	4524	17700
x"00",	-- Hex Addr	4525	17701
x"00",	-- Hex Addr	4526	17702
x"00",	-- Hex Addr	4527	17703
x"00",	-- Hex Addr	4528	17704
x"00",	-- Hex Addr	4529	17705
x"00",	-- Hex Addr	452A	17706
x"00",	-- Hex Addr	452B	17707
x"00",	-- Hex Addr	452C	17708
x"00",	-- Hex Addr	452D	17709
x"00",	-- Hex Addr	452E	17710
x"00",	-- Hex Addr	452F	17711
x"00",	-- Hex Addr	4530	17712
x"00",	-- Hex Addr	4531	17713
x"00",	-- Hex Addr	4532	17714
x"00",	-- Hex Addr	4533	17715
x"00",	-- Hex Addr	4534	17716
x"00",	-- Hex Addr	4535	17717
x"00",	-- Hex Addr	4536	17718
x"00",	-- Hex Addr	4537	17719
x"00",	-- Hex Addr	4538	17720
x"00",	-- Hex Addr	4539	17721
x"00",	-- Hex Addr	453A	17722
x"00",	-- Hex Addr	453B	17723
x"00",	-- Hex Addr	453C	17724
x"00",	-- Hex Addr	453D	17725
x"00",	-- Hex Addr	453E	17726
x"00",	-- Hex Addr	453F	17727
x"00",	-- Hex Addr	4540	17728
x"00",	-- Hex Addr	4541	17729
x"00",	-- Hex Addr	4542	17730
x"00",	-- Hex Addr	4543	17731
x"00",	-- Hex Addr	4544	17732
x"00",	-- Hex Addr	4545	17733
x"00",	-- Hex Addr	4546	17734
x"00",	-- Hex Addr	4547	17735
x"00",	-- Hex Addr	4548	17736
x"00",	-- Hex Addr	4549	17737
x"00",	-- Hex Addr	454A	17738
x"00",	-- Hex Addr	454B	17739
x"00",	-- Hex Addr	454C	17740
x"00",	-- Hex Addr	454D	17741
x"00",	-- Hex Addr	454E	17742
x"00",	-- Hex Addr	454F	17743
x"00",	-- Hex Addr	4550	17744
x"00",	-- Hex Addr	4551	17745
x"00",	-- Hex Addr	4552	17746
x"00",	-- Hex Addr	4553	17747
x"00",	-- Hex Addr	4554	17748
x"00",	-- Hex Addr	4555	17749
x"00",	-- Hex Addr	4556	17750
x"00",	-- Hex Addr	4557	17751
x"00",	-- Hex Addr	4558	17752
x"00",	-- Hex Addr	4559	17753
x"00",	-- Hex Addr	455A	17754
x"00",	-- Hex Addr	455B	17755
x"00",	-- Hex Addr	455C	17756
x"00",	-- Hex Addr	455D	17757
x"00",	-- Hex Addr	455E	17758
x"00",	-- Hex Addr	455F	17759
x"00",	-- Hex Addr	4560	17760
x"00",	-- Hex Addr	4561	17761
x"00",	-- Hex Addr	4562	17762
x"00",	-- Hex Addr	4563	17763
x"00",	-- Hex Addr	4564	17764
x"00",	-- Hex Addr	4565	17765
x"00",	-- Hex Addr	4566	17766
x"00",	-- Hex Addr	4567	17767
x"00",	-- Hex Addr	4568	17768
x"00",	-- Hex Addr	4569	17769
x"00",	-- Hex Addr	456A	17770
x"00",	-- Hex Addr	456B	17771
x"00",	-- Hex Addr	456C	17772
x"00",	-- Hex Addr	456D	17773
x"00",	-- Hex Addr	456E	17774
x"00",	-- Hex Addr	456F	17775
x"00",	-- Hex Addr	4570	17776
x"00",	-- Hex Addr	4571	17777
x"00",	-- Hex Addr	4572	17778
x"00",	-- Hex Addr	4573	17779
x"00",	-- Hex Addr	4574	17780
x"00",	-- Hex Addr	4575	17781
x"00",	-- Hex Addr	4576	17782
x"00",	-- Hex Addr	4577	17783
x"00",	-- Hex Addr	4578	17784
x"00",	-- Hex Addr	4579	17785
x"00",	-- Hex Addr	457A	17786
x"00",	-- Hex Addr	457B	17787
x"00",	-- Hex Addr	457C	17788
x"00",	-- Hex Addr	457D	17789
x"00",	-- Hex Addr	457E	17790
x"00",	-- Hex Addr	457F	17791
x"00",	-- Hex Addr	4580	17792
x"00",	-- Hex Addr	4581	17793
x"00",	-- Hex Addr	4582	17794
x"00",	-- Hex Addr	4583	17795
x"00",	-- Hex Addr	4584	17796
x"00",	-- Hex Addr	4585	17797
x"00",	-- Hex Addr	4586	17798
x"00",	-- Hex Addr	4587	17799
x"00",	-- Hex Addr	4588	17800
x"00",	-- Hex Addr	4589	17801
x"00",	-- Hex Addr	458A	17802
x"00",	-- Hex Addr	458B	17803
x"00",	-- Hex Addr	458C	17804
x"00",	-- Hex Addr	458D	17805
x"00",	-- Hex Addr	458E	17806
x"00",	-- Hex Addr	458F	17807
x"00",	-- Hex Addr	4590	17808
x"00",	-- Hex Addr	4591	17809
x"00",	-- Hex Addr	4592	17810
x"00",	-- Hex Addr	4593	17811
x"00",	-- Hex Addr	4594	17812
x"00",	-- Hex Addr	4595	17813
x"00",	-- Hex Addr	4596	17814
x"00",	-- Hex Addr	4597	17815
x"00",	-- Hex Addr	4598	17816
x"00",	-- Hex Addr	4599	17817
x"00",	-- Hex Addr	459A	17818
x"00",	-- Hex Addr	459B	17819
x"00",	-- Hex Addr	459C	17820
x"00",	-- Hex Addr	459D	17821
x"00",	-- Hex Addr	459E	17822
x"00",	-- Hex Addr	459F	17823
x"00",	-- Hex Addr	45A0	17824
x"00",	-- Hex Addr	45A1	17825
x"00",	-- Hex Addr	45A2	17826
x"00",	-- Hex Addr	45A3	17827
x"00",	-- Hex Addr	45A4	17828
x"00",	-- Hex Addr	45A5	17829
x"00",	-- Hex Addr	45A6	17830
x"00",	-- Hex Addr	45A7	17831
x"00",	-- Hex Addr	45A8	17832
x"00",	-- Hex Addr	45A9	17833
x"00",	-- Hex Addr	45AA	17834
x"00",	-- Hex Addr	45AB	17835
x"00",	-- Hex Addr	45AC	17836
x"00",	-- Hex Addr	45AD	17837
x"00",	-- Hex Addr	45AE	17838
x"00",	-- Hex Addr	45AF	17839
x"00",	-- Hex Addr	45B0	17840
x"00",	-- Hex Addr	45B1	17841
x"00",	-- Hex Addr	45B2	17842
x"00",	-- Hex Addr	45B3	17843
x"00",	-- Hex Addr	45B4	17844
x"00",	-- Hex Addr	45B5	17845
x"00",	-- Hex Addr	45B6	17846
x"00",	-- Hex Addr	45B7	17847
x"00",	-- Hex Addr	45B8	17848
x"00",	-- Hex Addr	45B9	17849
x"00",	-- Hex Addr	45BA	17850
x"00",	-- Hex Addr	45BB	17851
x"00",	-- Hex Addr	45BC	17852
x"00",	-- Hex Addr	45BD	17853
x"00",	-- Hex Addr	45BE	17854
x"00",	-- Hex Addr	45BF	17855
x"00",	-- Hex Addr	45C0	17856
x"00",	-- Hex Addr	45C1	17857
x"00",	-- Hex Addr	45C2	17858
x"00",	-- Hex Addr	45C3	17859
x"00",	-- Hex Addr	45C4	17860
x"00",	-- Hex Addr	45C5	17861
x"00",	-- Hex Addr	45C6	17862
x"00",	-- Hex Addr	45C7	17863
x"00",	-- Hex Addr	45C8	17864
x"00",	-- Hex Addr	45C9	17865
x"00",	-- Hex Addr	45CA	17866
x"00",	-- Hex Addr	45CB	17867
x"00",	-- Hex Addr	45CC	17868
x"00",	-- Hex Addr	45CD	17869
x"00",	-- Hex Addr	45CE	17870
x"00",	-- Hex Addr	45CF	17871
x"00",	-- Hex Addr	45D0	17872
x"00",	-- Hex Addr	45D1	17873
x"00",	-- Hex Addr	45D2	17874
x"00",	-- Hex Addr	45D3	17875
x"00",	-- Hex Addr	45D4	17876
x"00",	-- Hex Addr	45D5	17877
x"00",	-- Hex Addr	45D6	17878
x"00",	-- Hex Addr	45D7	17879
x"00",	-- Hex Addr	45D8	17880
x"00",	-- Hex Addr	45D9	17881
x"00",	-- Hex Addr	45DA	17882
x"00",	-- Hex Addr	45DB	17883
x"00",	-- Hex Addr	45DC	17884
x"00",	-- Hex Addr	45DD	17885
x"00",	-- Hex Addr	45DE	17886
x"00",	-- Hex Addr	45DF	17887
x"00",	-- Hex Addr	45E0	17888
x"00",	-- Hex Addr	45E1	17889
x"00",	-- Hex Addr	45E2	17890
x"00",	-- Hex Addr	45E3	17891
x"00",	-- Hex Addr	45E4	17892
x"00",	-- Hex Addr	45E5	17893
x"00",	-- Hex Addr	45E6	17894
x"00",	-- Hex Addr	45E7	17895
x"00",	-- Hex Addr	45E8	17896
x"00",	-- Hex Addr	45E9	17897
x"00",	-- Hex Addr	45EA	17898
x"00",	-- Hex Addr	45EB	17899
x"00",	-- Hex Addr	45EC	17900
x"00",	-- Hex Addr	45ED	17901
x"00",	-- Hex Addr	45EE	17902
x"00",	-- Hex Addr	45EF	17903
x"00",	-- Hex Addr	45F0	17904
x"00",	-- Hex Addr	45F1	17905
x"00",	-- Hex Addr	45F2	17906
x"00",	-- Hex Addr	45F3	17907
x"00",	-- Hex Addr	45F4	17908
x"00",	-- Hex Addr	45F5	17909
x"00",	-- Hex Addr	45F6	17910
x"00",	-- Hex Addr	45F7	17911
x"00",	-- Hex Addr	45F8	17912
x"00",	-- Hex Addr	45F9	17913
x"00",	-- Hex Addr	45FA	17914
x"00",	-- Hex Addr	45FB	17915
x"00",	-- Hex Addr	45FC	17916
x"00",	-- Hex Addr	45FD	17917
x"00",	-- Hex Addr	45FE	17918
x"00",	-- Hex Addr	45FF	17919
x"00",	-- Hex Addr	4600	17920
x"00",	-- Hex Addr	4601	17921
x"00",	-- Hex Addr	4602	17922
x"00",	-- Hex Addr	4603	17923
x"00",	-- Hex Addr	4604	17924
x"00",	-- Hex Addr	4605	17925
x"00",	-- Hex Addr	4606	17926
x"00",	-- Hex Addr	4607	17927
x"00",	-- Hex Addr	4608	17928
x"00",	-- Hex Addr	4609	17929
x"00",	-- Hex Addr	460A	17930
x"00",	-- Hex Addr	460B	17931
x"00",	-- Hex Addr	460C	17932
x"00",	-- Hex Addr	460D	17933
x"00",	-- Hex Addr	460E	17934
x"00",	-- Hex Addr	460F	17935
x"00",	-- Hex Addr	4610	17936
x"00",	-- Hex Addr	4611	17937
x"00",	-- Hex Addr	4612	17938
x"00",	-- Hex Addr	4613	17939
x"00",	-- Hex Addr	4614	17940
x"00",	-- Hex Addr	4615	17941
x"00",	-- Hex Addr	4616	17942
x"00",	-- Hex Addr	4617	17943
x"00",	-- Hex Addr	4618	17944
x"00",	-- Hex Addr	4619	17945
x"00",	-- Hex Addr	461A	17946
x"00",	-- Hex Addr	461B	17947
x"00",	-- Hex Addr	461C	17948
x"00",	-- Hex Addr	461D	17949
x"00",	-- Hex Addr	461E	17950
x"00",	-- Hex Addr	461F	17951
x"00",	-- Hex Addr	4620	17952
x"00",	-- Hex Addr	4621	17953
x"00",	-- Hex Addr	4622	17954
x"00",	-- Hex Addr	4623	17955
x"00",	-- Hex Addr	4624	17956
x"00",	-- Hex Addr	4625	17957
x"00",	-- Hex Addr	4626	17958
x"00",	-- Hex Addr	4627	17959
x"00",	-- Hex Addr	4628	17960
x"00",	-- Hex Addr	4629	17961
x"00",	-- Hex Addr	462A	17962
x"00",	-- Hex Addr	462B	17963
x"00",	-- Hex Addr	462C	17964
x"00",	-- Hex Addr	462D	17965
x"00",	-- Hex Addr	462E	17966
x"00",	-- Hex Addr	462F	17967
x"00",	-- Hex Addr	4630	17968
x"00",	-- Hex Addr	4631	17969
x"00",	-- Hex Addr	4632	17970
x"00",	-- Hex Addr	4633	17971
x"00",	-- Hex Addr	4634	17972
x"00",	-- Hex Addr	4635	17973
x"00",	-- Hex Addr	4636	17974
x"00",	-- Hex Addr	4637	17975
x"00",	-- Hex Addr	4638	17976
x"00",	-- Hex Addr	4639	17977
x"00",	-- Hex Addr	463A	17978
x"00",	-- Hex Addr	463B	17979
x"00",	-- Hex Addr	463C	17980
x"00",	-- Hex Addr	463D	17981
x"00",	-- Hex Addr	463E	17982
x"00",	-- Hex Addr	463F	17983
x"00",	-- Hex Addr	4640	17984
x"00",	-- Hex Addr	4641	17985
x"00",	-- Hex Addr	4642	17986
x"00",	-- Hex Addr	4643	17987
x"00",	-- Hex Addr	4644	17988
x"00",	-- Hex Addr	4645	17989
x"00",	-- Hex Addr	4646	17990
x"00",	-- Hex Addr	4647	17991
x"00",	-- Hex Addr	4648	17992
x"00",	-- Hex Addr	4649	17993
x"00",	-- Hex Addr	464A	17994
x"00",	-- Hex Addr	464B	17995
x"00",	-- Hex Addr	464C	17996
x"00",	-- Hex Addr	464D	17997
x"00",	-- Hex Addr	464E	17998
x"00",	-- Hex Addr	464F	17999
x"00",	-- Hex Addr	4650	18000
x"00",	-- Hex Addr	4651	18001
x"00",	-- Hex Addr	4652	18002
x"00",	-- Hex Addr	4653	18003
x"00",	-- Hex Addr	4654	18004
x"00",	-- Hex Addr	4655	18005
x"00",	-- Hex Addr	4656	18006
x"00",	-- Hex Addr	4657	18007
x"00",	-- Hex Addr	4658	18008
x"00",	-- Hex Addr	4659	18009
x"00",	-- Hex Addr	465A	18010
x"00",	-- Hex Addr	465B	18011
x"00",	-- Hex Addr	465C	18012
x"00",	-- Hex Addr	465D	18013
x"00",	-- Hex Addr	465E	18014
x"00",	-- Hex Addr	465F	18015
x"00",	-- Hex Addr	4660	18016
x"00",	-- Hex Addr	4661	18017
x"00",	-- Hex Addr	4662	18018
x"00",	-- Hex Addr	4663	18019
x"00",	-- Hex Addr	4664	18020
x"00",	-- Hex Addr	4665	18021
x"00",	-- Hex Addr	4666	18022
x"00",	-- Hex Addr	4667	18023
x"00",	-- Hex Addr	4668	18024
x"00",	-- Hex Addr	4669	18025
x"00",	-- Hex Addr	466A	18026
x"00",	-- Hex Addr	466B	18027
x"00",	-- Hex Addr	466C	18028
x"00",	-- Hex Addr	466D	18029
x"00",	-- Hex Addr	466E	18030
x"00",	-- Hex Addr	466F	18031
x"00",	-- Hex Addr	4670	18032
x"00",	-- Hex Addr	4671	18033
x"00",	-- Hex Addr	4672	18034
x"00",	-- Hex Addr	4673	18035
x"00",	-- Hex Addr	4674	18036
x"00",	-- Hex Addr	4675	18037
x"00",	-- Hex Addr	4676	18038
x"00",	-- Hex Addr	4677	18039
x"00",	-- Hex Addr	4678	18040
x"00",	-- Hex Addr	4679	18041
x"00",	-- Hex Addr	467A	18042
x"00",	-- Hex Addr	467B	18043
x"00",	-- Hex Addr	467C	18044
x"00",	-- Hex Addr	467D	18045
x"00",	-- Hex Addr	467E	18046
x"00",	-- Hex Addr	467F	18047
x"00",	-- Hex Addr	4680	18048
x"00",	-- Hex Addr	4681	18049
x"00",	-- Hex Addr	4682	18050
x"00",	-- Hex Addr	4683	18051
x"00",	-- Hex Addr	4684	18052
x"00",	-- Hex Addr	4685	18053
x"00",	-- Hex Addr	4686	18054
x"00",	-- Hex Addr	4687	18055
x"00",	-- Hex Addr	4688	18056
x"00",	-- Hex Addr	4689	18057
x"00",	-- Hex Addr	468A	18058
x"00",	-- Hex Addr	468B	18059
x"00",	-- Hex Addr	468C	18060
x"00",	-- Hex Addr	468D	18061
x"00",	-- Hex Addr	468E	18062
x"00",	-- Hex Addr	468F	18063
x"00",	-- Hex Addr	4690	18064
x"00",	-- Hex Addr	4691	18065
x"00",	-- Hex Addr	4692	18066
x"00",	-- Hex Addr	4693	18067
x"00",	-- Hex Addr	4694	18068
x"00",	-- Hex Addr	4695	18069
x"00",	-- Hex Addr	4696	18070
x"00",	-- Hex Addr	4697	18071
x"00",	-- Hex Addr	4698	18072
x"00",	-- Hex Addr	4699	18073
x"00",	-- Hex Addr	469A	18074
x"00",	-- Hex Addr	469B	18075
x"00",	-- Hex Addr	469C	18076
x"00",	-- Hex Addr	469D	18077
x"00",	-- Hex Addr	469E	18078
x"00",	-- Hex Addr	469F	18079
x"00",	-- Hex Addr	46A0	18080
x"00",	-- Hex Addr	46A1	18081
x"00",	-- Hex Addr	46A2	18082
x"00",	-- Hex Addr	46A3	18083
x"00",	-- Hex Addr	46A4	18084
x"00",	-- Hex Addr	46A5	18085
x"00",	-- Hex Addr	46A6	18086
x"00",	-- Hex Addr	46A7	18087
x"00",	-- Hex Addr	46A8	18088
x"00",	-- Hex Addr	46A9	18089
x"00",	-- Hex Addr	46AA	18090
x"00",	-- Hex Addr	46AB	18091
x"00",	-- Hex Addr	46AC	18092
x"00",	-- Hex Addr	46AD	18093
x"00",	-- Hex Addr	46AE	18094
x"00",	-- Hex Addr	46AF	18095
x"00",	-- Hex Addr	46B0	18096
x"00",	-- Hex Addr	46B1	18097
x"00",	-- Hex Addr	46B2	18098
x"00",	-- Hex Addr	46B3	18099
x"00",	-- Hex Addr	46B4	18100
x"00",	-- Hex Addr	46B5	18101
x"00",	-- Hex Addr	46B6	18102
x"00",	-- Hex Addr	46B7	18103
x"00",	-- Hex Addr	46B8	18104
x"00",	-- Hex Addr	46B9	18105
x"00",	-- Hex Addr	46BA	18106
x"00",	-- Hex Addr	46BB	18107
x"00",	-- Hex Addr	46BC	18108
x"00",	-- Hex Addr	46BD	18109
x"00",	-- Hex Addr	46BE	18110
x"00",	-- Hex Addr	46BF	18111
x"00",	-- Hex Addr	46C0	18112
x"00",	-- Hex Addr	46C1	18113
x"00",	-- Hex Addr	46C2	18114
x"00",	-- Hex Addr	46C3	18115
x"00",	-- Hex Addr	46C4	18116
x"00",	-- Hex Addr	46C5	18117
x"00",	-- Hex Addr	46C6	18118
x"00",	-- Hex Addr	46C7	18119
x"00",	-- Hex Addr	46C8	18120
x"00",	-- Hex Addr	46C9	18121
x"00",	-- Hex Addr	46CA	18122
x"00",	-- Hex Addr	46CB	18123
x"00",	-- Hex Addr	46CC	18124
x"00",	-- Hex Addr	46CD	18125
x"00",	-- Hex Addr	46CE	18126
x"00",	-- Hex Addr	46CF	18127
x"00",	-- Hex Addr	46D0	18128
x"00",	-- Hex Addr	46D1	18129
x"00",	-- Hex Addr	46D2	18130
x"00",	-- Hex Addr	46D3	18131
x"00",	-- Hex Addr	46D4	18132
x"00",	-- Hex Addr	46D5	18133
x"00",	-- Hex Addr	46D6	18134
x"00",	-- Hex Addr	46D7	18135
x"00",	-- Hex Addr	46D8	18136
x"00",	-- Hex Addr	46D9	18137
x"00",	-- Hex Addr	46DA	18138
x"00",	-- Hex Addr	46DB	18139
x"00",	-- Hex Addr	46DC	18140
x"00",	-- Hex Addr	46DD	18141
x"00",	-- Hex Addr	46DE	18142
x"00",	-- Hex Addr	46DF	18143
x"00",	-- Hex Addr	46E0	18144
x"00",	-- Hex Addr	46E1	18145
x"00",	-- Hex Addr	46E2	18146
x"00",	-- Hex Addr	46E3	18147
x"00",	-- Hex Addr	46E4	18148
x"00",	-- Hex Addr	46E5	18149
x"00",	-- Hex Addr	46E6	18150
x"00",	-- Hex Addr	46E7	18151
x"00",	-- Hex Addr	46E8	18152
x"00",	-- Hex Addr	46E9	18153
x"00",	-- Hex Addr	46EA	18154
x"00",	-- Hex Addr	46EB	18155
x"00",	-- Hex Addr	46EC	18156
x"00",	-- Hex Addr	46ED	18157
x"00",	-- Hex Addr	46EE	18158
x"00",	-- Hex Addr	46EF	18159
x"00",	-- Hex Addr	46F0	18160
x"00",	-- Hex Addr	46F1	18161
x"00",	-- Hex Addr	46F2	18162
x"00",	-- Hex Addr	46F3	18163
x"00",	-- Hex Addr	46F4	18164
x"00",	-- Hex Addr	46F5	18165
x"00",	-- Hex Addr	46F6	18166
x"00",	-- Hex Addr	46F7	18167
x"00",	-- Hex Addr	46F8	18168
x"00",	-- Hex Addr	46F9	18169
x"00",	-- Hex Addr	46FA	18170
x"00",	-- Hex Addr	46FB	18171
x"00",	-- Hex Addr	46FC	18172
x"00",	-- Hex Addr	46FD	18173
x"00",	-- Hex Addr	46FE	18174
x"00",	-- Hex Addr	46FF	18175
x"00",	-- Hex Addr	4700	18176
x"00",	-- Hex Addr	4701	18177
x"00",	-- Hex Addr	4702	18178
x"00",	-- Hex Addr	4703	18179
x"00",	-- Hex Addr	4704	18180
x"00",	-- Hex Addr	4705	18181
x"00",	-- Hex Addr	4706	18182
x"00",	-- Hex Addr	4707	18183
x"00",	-- Hex Addr	4708	18184
x"00",	-- Hex Addr	4709	18185
x"00",	-- Hex Addr	470A	18186
x"00",	-- Hex Addr	470B	18187
x"00",	-- Hex Addr	470C	18188
x"00",	-- Hex Addr	470D	18189
x"00",	-- Hex Addr	470E	18190
x"00",	-- Hex Addr	470F	18191
x"00",	-- Hex Addr	4710	18192
x"00",	-- Hex Addr	4711	18193
x"00",	-- Hex Addr	4712	18194
x"00",	-- Hex Addr	4713	18195
x"00",	-- Hex Addr	4714	18196
x"00",	-- Hex Addr	4715	18197
x"00",	-- Hex Addr	4716	18198
x"00",	-- Hex Addr	4717	18199
x"00",	-- Hex Addr	4718	18200
x"00",	-- Hex Addr	4719	18201
x"00",	-- Hex Addr	471A	18202
x"00",	-- Hex Addr	471B	18203
x"00",	-- Hex Addr	471C	18204
x"00",	-- Hex Addr	471D	18205
x"00",	-- Hex Addr	471E	18206
x"00",	-- Hex Addr	471F	18207
x"00",	-- Hex Addr	4720	18208
x"00",	-- Hex Addr	4721	18209
x"00",	-- Hex Addr	4722	18210
x"00",	-- Hex Addr	4723	18211
x"00",	-- Hex Addr	4724	18212
x"00",	-- Hex Addr	4725	18213
x"00",	-- Hex Addr	4726	18214
x"00",	-- Hex Addr	4727	18215
x"00",	-- Hex Addr	4728	18216
x"00",	-- Hex Addr	4729	18217
x"00",	-- Hex Addr	472A	18218
x"00",	-- Hex Addr	472B	18219
x"00",	-- Hex Addr	472C	18220
x"00",	-- Hex Addr	472D	18221
x"00",	-- Hex Addr	472E	18222
x"00",	-- Hex Addr	472F	18223
x"00",	-- Hex Addr	4730	18224
x"00",	-- Hex Addr	4731	18225
x"00",	-- Hex Addr	4732	18226
x"00",	-- Hex Addr	4733	18227
x"00",	-- Hex Addr	4734	18228
x"00",	-- Hex Addr	4735	18229
x"00",	-- Hex Addr	4736	18230
x"00",	-- Hex Addr	4737	18231
x"00",	-- Hex Addr	4738	18232
x"00",	-- Hex Addr	4739	18233
x"00",	-- Hex Addr	473A	18234
x"00",	-- Hex Addr	473B	18235
x"00",	-- Hex Addr	473C	18236
x"00",	-- Hex Addr	473D	18237
x"00",	-- Hex Addr	473E	18238
x"00",	-- Hex Addr	473F	18239
x"00",	-- Hex Addr	4740	18240
x"00",	-- Hex Addr	4741	18241
x"00",	-- Hex Addr	4742	18242
x"00",	-- Hex Addr	4743	18243
x"00",	-- Hex Addr	4744	18244
x"00",	-- Hex Addr	4745	18245
x"00",	-- Hex Addr	4746	18246
x"00",	-- Hex Addr	4747	18247
x"00",	-- Hex Addr	4748	18248
x"00",	-- Hex Addr	4749	18249
x"00",	-- Hex Addr	474A	18250
x"00",	-- Hex Addr	474B	18251
x"00",	-- Hex Addr	474C	18252
x"00",	-- Hex Addr	474D	18253
x"00",	-- Hex Addr	474E	18254
x"00",	-- Hex Addr	474F	18255
x"00",	-- Hex Addr	4750	18256
x"00",	-- Hex Addr	4751	18257
x"00",	-- Hex Addr	4752	18258
x"00",	-- Hex Addr	4753	18259
x"00",	-- Hex Addr	4754	18260
x"00",	-- Hex Addr	4755	18261
x"00",	-- Hex Addr	4756	18262
x"00",	-- Hex Addr	4757	18263
x"00",	-- Hex Addr	4758	18264
x"00",	-- Hex Addr	4759	18265
x"00",	-- Hex Addr	475A	18266
x"00",	-- Hex Addr	475B	18267
x"00",	-- Hex Addr	475C	18268
x"00",	-- Hex Addr	475D	18269
x"00",	-- Hex Addr	475E	18270
x"00",	-- Hex Addr	475F	18271
x"00",	-- Hex Addr	4760	18272
x"00",	-- Hex Addr	4761	18273
x"00",	-- Hex Addr	4762	18274
x"00",	-- Hex Addr	4763	18275
x"00",	-- Hex Addr	4764	18276
x"00",	-- Hex Addr	4765	18277
x"00",	-- Hex Addr	4766	18278
x"00",	-- Hex Addr	4767	18279
x"00",	-- Hex Addr	4768	18280
x"00",	-- Hex Addr	4769	18281
x"00",	-- Hex Addr	476A	18282
x"00",	-- Hex Addr	476B	18283
x"00",	-- Hex Addr	476C	18284
x"00",	-- Hex Addr	476D	18285
x"00",	-- Hex Addr	476E	18286
x"00",	-- Hex Addr	476F	18287
x"00",	-- Hex Addr	4770	18288
x"00",	-- Hex Addr	4771	18289
x"00",	-- Hex Addr	4772	18290
x"00",	-- Hex Addr	4773	18291
x"00",	-- Hex Addr	4774	18292
x"00",	-- Hex Addr	4775	18293
x"00",	-- Hex Addr	4776	18294
x"00",	-- Hex Addr	4777	18295
x"00",	-- Hex Addr	4778	18296
x"00",	-- Hex Addr	4779	18297
x"00",	-- Hex Addr	477A	18298
x"00",	-- Hex Addr	477B	18299
x"00",	-- Hex Addr	477C	18300
x"00",	-- Hex Addr	477D	18301
x"00",	-- Hex Addr	477E	18302
x"00",	-- Hex Addr	477F	18303
x"00",	-- Hex Addr	4780	18304
x"00",	-- Hex Addr	4781	18305
x"00",	-- Hex Addr	4782	18306
x"00",	-- Hex Addr	4783	18307
x"00",	-- Hex Addr	4784	18308
x"00",	-- Hex Addr	4785	18309
x"00",	-- Hex Addr	4786	18310
x"00",	-- Hex Addr	4787	18311
x"00",	-- Hex Addr	4788	18312
x"00",	-- Hex Addr	4789	18313
x"00",	-- Hex Addr	478A	18314
x"00",	-- Hex Addr	478B	18315
x"00",	-- Hex Addr	478C	18316
x"00",	-- Hex Addr	478D	18317
x"00",	-- Hex Addr	478E	18318
x"00",	-- Hex Addr	478F	18319
x"00",	-- Hex Addr	4790	18320
x"00",	-- Hex Addr	4791	18321
x"00",	-- Hex Addr	4792	18322
x"00",	-- Hex Addr	4793	18323
x"00",	-- Hex Addr	4794	18324
x"00",	-- Hex Addr	4795	18325
x"00",	-- Hex Addr	4796	18326
x"00",	-- Hex Addr	4797	18327
x"00",	-- Hex Addr	4798	18328
x"00",	-- Hex Addr	4799	18329
x"00",	-- Hex Addr	479A	18330
x"00",	-- Hex Addr	479B	18331
x"00",	-- Hex Addr	479C	18332
x"00",	-- Hex Addr	479D	18333
x"00",	-- Hex Addr	479E	18334
x"00",	-- Hex Addr	479F	18335
x"00",	-- Hex Addr	47A0	18336
x"00",	-- Hex Addr	47A1	18337
x"00",	-- Hex Addr	47A2	18338
x"00",	-- Hex Addr	47A3	18339
x"00",	-- Hex Addr	47A4	18340
x"00",	-- Hex Addr	47A5	18341
x"00",	-- Hex Addr	47A6	18342
x"00",	-- Hex Addr	47A7	18343
x"00",	-- Hex Addr	47A8	18344
x"00",	-- Hex Addr	47A9	18345
x"00",	-- Hex Addr	47AA	18346
x"00",	-- Hex Addr	47AB	18347
x"00",	-- Hex Addr	47AC	18348
x"00",	-- Hex Addr	47AD	18349
x"00",	-- Hex Addr	47AE	18350
x"00",	-- Hex Addr	47AF	18351
x"00",	-- Hex Addr	47B0	18352
x"00",	-- Hex Addr	47B1	18353
x"00",	-- Hex Addr	47B2	18354
x"00",	-- Hex Addr	47B3	18355
x"00",	-- Hex Addr	47B4	18356
x"00",	-- Hex Addr	47B5	18357
x"00",	-- Hex Addr	47B6	18358
x"00",	-- Hex Addr	47B7	18359
x"00",	-- Hex Addr	47B8	18360
x"00",	-- Hex Addr	47B9	18361
x"00",	-- Hex Addr	47BA	18362
x"00",	-- Hex Addr	47BB	18363
x"00",	-- Hex Addr	47BC	18364
x"00",	-- Hex Addr	47BD	18365
x"00",	-- Hex Addr	47BE	18366
x"00",	-- Hex Addr	47BF	18367
x"00",	-- Hex Addr	47C0	18368
x"00",	-- Hex Addr	47C1	18369
x"00",	-- Hex Addr	47C2	18370
x"00",	-- Hex Addr	47C3	18371
x"00",	-- Hex Addr	47C4	18372
x"00",	-- Hex Addr	47C5	18373
x"00",	-- Hex Addr	47C6	18374
x"00",	-- Hex Addr	47C7	18375
x"00",	-- Hex Addr	47C8	18376
x"00",	-- Hex Addr	47C9	18377
x"00",	-- Hex Addr	47CA	18378
x"00",	-- Hex Addr	47CB	18379
x"00",	-- Hex Addr	47CC	18380
x"00",	-- Hex Addr	47CD	18381
x"00",	-- Hex Addr	47CE	18382
x"00",	-- Hex Addr	47CF	18383
x"00",	-- Hex Addr	47D0	18384
x"00",	-- Hex Addr	47D1	18385
x"00",	-- Hex Addr	47D2	18386
x"00",	-- Hex Addr	47D3	18387
x"00",	-- Hex Addr	47D4	18388
x"00",	-- Hex Addr	47D5	18389
x"00",	-- Hex Addr	47D6	18390
x"00",	-- Hex Addr	47D7	18391
x"00",	-- Hex Addr	47D8	18392
x"00",	-- Hex Addr	47D9	18393
x"00",	-- Hex Addr	47DA	18394
x"00",	-- Hex Addr	47DB	18395
x"00",	-- Hex Addr	47DC	18396
x"00",	-- Hex Addr	47DD	18397
x"00",	-- Hex Addr	47DE	18398
x"00",	-- Hex Addr	47DF	18399
x"00",	-- Hex Addr	47E0	18400
x"00",	-- Hex Addr	47E1	18401
x"00",	-- Hex Addr	47E2	18402
x"00",	-- Hex Addr	47E3	18403
x"00",	-- Hex Addr	47E4	18404
x"00",	-- Hex Addr	47E5	18405
x"00",	-- Hex Addr	47E6	18406
x"00",	-- Hex Addr	47E7	18407
x"00",	-- Hex Addr	47E8	18408
x"00",	-- Hex Addr	47E9	18409
x"00",	-- Hex Addr	47EA	18410
x"00",	-- Hex Addr	47EB	18411
x"00",	-- Hex Addr	47EC	18412
x"00",	-- Hex Addr	47ED	18413
x"00",	-- Hex Addr	47EE	18414
x"00",	-- Hex Addr	47EF	18415
x"00",	-- Hex Addr	47F0	18416
x"00",	-- Hex Addr	47F1	18417
x"00",	-- Hex Addr	47F2	18418
x"00",	-- Hex Addr	47F3	18419
x"00",	-- Hex Addr	47F4	18420
x"00",	-- Hex Addr	47F5	18421
x"00",	-- Hex Addr	47F6	18422
x"00",	-- Hex Addr	47F7	18423
x"00",	-- Hex Addr	47F8	18424
x"00",	-- Hex Addr	47F9	18425
x"00",	-- Hex Addr	47FA	18426
x"00",	-- Hex Addr	47FB	18427
x"00",	-- Hex Addr	47FC	18428
x"00",	-- Hex Addr	47FD	18429
x"00",	-- Hex Addr	47FE	18430
x"00",	-- Hex Addr	47FF	18431
x"00",	-- Hex Addr	4800	18432
x"00",	-- Hex Addr	4801	18433
x"00",	-- Hex Addr	4802	18434
x"00",	-- Hex Addr	4803	18435
x"00",	-- Hex Addr	4804	18436
x"00",	-- Hex Addr	4805	18437
x"00",	-- Hex Addr	4806	18438
x"00",	-- Hex Addr	4807	18439
x"00",	-- Hex Addr	4808	18440
x"00",	-- Hex Addr	4809	18441
x"00",	-- Hex Addr	480A	18442
x"00",	-- Hex Addr	480B	18443
x"00",	-- Hex Addr	480C	18444
x"00",	-- Hex Addr	480D	18445
x"00",	-- Hex Addr	480E	18446
x"00",	-- Hex Addr	480F	18447
x"00",	-- Hex Addr	4810	18448
x"00",	-- Hex Addr	4811	18449
x"00",	-- Hex Addr	4812	18450
x"00",	-- Hex Addr	4813	18451
x"00",	-- Hex Addr	4814	18452
x"00",	-- Hex Addr	4815	18453
x"00",	-- Hex Addr	4816	18454
x"00",	-- Hex Addr	4817	18455
x"00",	-- Hex Addr	4818	18456
x"00",	-- Hex Addr	4819	18457
x"00",	-- Hex Addr	481A	18458
x"00",	-- Hex Addr	481B	18459
x"00",	-- Hex Addr	481C	18460
x"00",	-- Hex Addr	481D	18461
x"00",	-- Hex Addr	481E	18462
x"00",	-- Hex Addr	481F	18463
x"00",	-- Hex Addr	4820	18464
x"00",	-- Hex Addr	4821	18465
x"00",	-- Hex Addr	4822	18466
x"00",	-- Hex Addr	4823	18467
x"00",	-- Hex Addr	4824	18468
x"00",	-- Hex Addr	4825	18469
x"00",	-- Hex Addr	4826	18470
x"00",	-- Hex Addr	4827	18471
x"00",	-- Hex Addr	4828	18472
x"00",	-- Hex Addr	4829	18473
x"00",	-- Hex Addr	482A	18474
x"00",	-- Hex Addr	482B	18475
x"00",	-- Hex Addr	482C	18476
x"00",	-- Hex Addr	482D	18477
x"00",	-- Hex Addr	482E	18478
x"00",	-- Hex Addr	482F	18479
x"00",	-- Hex Addr	4830	18480
x"00",	-- Hex Addr	4831	18481
x"00",	-- Hex Addr	4832	18482
x"00",	-- Hex Addr	4833	18483
x"00",	-- Hex Addr	4834	18484
x"00",	-- Hex Addr	4835	18485
x"00",	-- Hex Addr	4836	18486
x"00",	-- Hex Addr	4837	18487
x"00",	-- Hex Addr	4838	18488
x"00",	-- Hex Addr	4839	18489
x"00",	-- Hex Addr	483A	18490
x"00",	-- Hex Addr	483B	18491
x"00",	-- Hex Addr	483C	18492
x"00",	-- Hex Addr	483D	18493
x"00",	-- Hex Addr	483E	18494
x"00",	-- Hex Addr	483F	18495
x"00",	-- Hex Addr	4840	18496
x"00",	-- Hex Addr	4841	18497
x"00",	-- Hex Addr	4842	18498
x"00",	-- Hex Addr	4843	18499
x"00",	-- Hex Addr	4844	18500
x"00",	-- Hex Addr	4845	18501
x"00",	-- Hex Addr	4846	18502
x"00",	-- Hex Addr	4847	18503
x"00",	-- Hex Addr	4848	18504
x"00",	-- Hex Addr	4849	18505
x"00",	-- Hex Addr	484A	18506
x"00",	-- Hex Addr	484B	18507
x"00",	-- Hex Addr	484C	18508
x"00",	-- Hex Addr	484D	18509
x"00",	-- Hex Addr	484E	18510
x"00",	-- Hex Addr	484F	18511
x"00",	-- Hex Addr	4850	18512
x"00",	-- Hex Addr	4851	18513
x"00",	-- Hex Addr	4852	18514
x"00",	-- Hex Addr	4853	18515
x"00",	-- Hex Addr	4854	18516
x"00",	-- Hex Addr	4855	18517
x"00",	-- Hex Addr	4856	18518
x"00",	-- Hex Addr	4857	18519
x"00",	-- Hex Addr	4858	18520
x"00",	-- Hex Addr	4859	18521
x"00",	-- Hex Addr	485A	18522
x"00",	-- Hex Addr	485B	18523
x"00",	-- Hex Addr	485C	18524
x"00",	-- Hex Addr	485D	18525
x"00",	-- Hex Addr	485E	18526
x"00",	-- Hex Addr	485F	18527
x"00",	-- Hex Addr	4860	18528
x"00",	-- Hex Addr	4861	18529
x"00",	-- Hex Addr	4862	18530
x"00",	-- Hex Addr	4863	18531
x"00",	-- Hex Addr	4864	18532
x"00",	-- Hex Addr	4865	18533
x"00",	-- Hex Addr	4866	18534
x"00",	-- Hex Addr	4867	18535
x"00",	-- Hex Addr	4868	18536
x"00",	-- Hex Addr	4869	18537
x"00",	-- Hex Addr	486A	18538
x"00",	-- Hex Addr	486B	18539
x"00",	-- Hex Addr	486C	18540
x"00",	-- Hex Addr	486D	18541
x"00",	-- Hex Addr	486E	18542
x"00",	-- Hex Addr	486F	18543
x"00",	-- Hex Addr	4870	18544
x"00",	-- Hex Addr	4871	18545
x"00",	-- Hex Addr	4872	18546
x"00",	-- Hex Addr	4873	18547
x"00",	-- Hex Addr	4874	18548
x"00",	-- Hex Addr	4875	18549
x"00",	-- Hex Addr	4876	18550
x"00",	-- Hex Addr	4877	18551
x"00",	-- Hex Addr	4878	18552
x"00",	-- Hex Addr	4879	18553
x"00",	-- Hex Addr	487A	18554
x"00",	-- Hex Addr	487B	18555
x"00",	-- Hex Addr	487C	18556
x"00",	-- Hex Addr	487D	18557
x"00",	-- Hex Addr	487E	18558
x"00",	-- Hex Addr	487F	18559
x"00",	-- Hex Addr	4880	18560
x"00",	-- Hex Addr	4881	18561
x"00",	-- Hex Addr	4882	18562
x"00",	-- Hex Addr	4883	18563
x"00",	-- Hex Addr	4884	18564
x"00",	-- Hex Addr	4885	18565
x"00",	-- Hex Addr	4886	18566
x"00",	-- Hex Addr	4887	18567
x"00",	-- Hex Addr	4888	18568
x"00",	-- Hex Addr	4889	18569
x"00",	-- Hex Addr	488A	18570
x"00",	-- Hex Addr	488B	18571
x"00",	-- Hex Addr	488C	18572
x"00",	-- Hex Addr	488D	18573
x"00",	-- Hex Addr	488E	18574
x"00",	-- Hex Addr	488F	18575
x"00",	-- Hex Addr	4890	18576
x"00",	-- Hex Addr	4891	18577
x"00",	-- Hex Addr	4892	18578
x"00",	-- Hex Addr	4893	18579
x"00",	-- Hex Addr	4894	18580
x"00",	-- Hex Addr	4895	18581
x"00",	-- Hex Addr	4896	18582
x"00",	-- Hex Addr	4897	18583
x"00",	-- Hex Addr	4898	18584
x"00",	-- Hex Addr	4899	18585
x"00",	-- Hex Addr	489A	18586
x"00",	-- Hex Addr	489B	18587
x"00",	-- Hex Addr	489C	18588
x"00",	-- Hex Addr	489D	18589
x"00",	-- Hex Addr	489E	18590
x"00",	-- Hex Addr	489F	18591
x"00",	-- Hex Addr	48A0	18592
x"00",	-- Hex Addr	48A1	18593
x"00",	-- Hex Addr	48A2	18594
x"00",	-- Hex Addr	48A3	18595
x"00",	-- Hex Addr	48A4	18596
x"00",	-- Hex Addr	48A5	18597
x"00",	-- Hex Addr	48A6	18598
x"00",	-- Hex Addr	48A7	18599
x"00",	-- Hex Addr	48A8	18600
x"00",	-- Hex Addr	48A9	18601
x"00",	-- Hex Addr	48AA	18602
x"00",	-- Hex Addr	48AB	18603
x"00",	-- Hex Addr	48AC	18604
x"00",	-- Hex Addr	48AD	18605
x"00",	-- Hex Addr	48AE	18606
x"00",	-- Hex Addr	48AF	18607
x"00",	-- Hex Addr	48B0	18608
x"00",	-- Hex Addr	48B1	18609
x"00",	-- Hex Addr	48B2	18610
x"00",	-- Hex Addr	48B3	18611
x"00",	-- Hex Addr	48B4	18612
x"00",	-- Hex Addr	48B5	18613
x"00",	-- Hex Addr	48B6	18614
x"00",	-- Hex Addr	48B7	18615
x"00",	-- Hex Addr	48B8	18616
x"00",	-- Hex Addr	48B9	18617
x"00",	-- Hex Addr	48BA	18618
x"00",	-- Hex Addr	48BB	18619
x"00",	-- Hex Addr	48BC	18620
x"00",	-- Hex Addr	48BD	18621
x"00",	-- Hex Addr	48BE	18622
x"00",	-- Hex Addr	48BF	18623
x"00",	-- Hex Addr	48C0	18624
x"00",	-- Hex Addr	48C1	18625
x"00",	-- Hex Addr	48C2	18626
x"00",	-- Hex Addr	48C3	18627
x"00",	-- Hex Addr	48C4	18628
x"00",	-- Hex Addr	48C5	18629
x"00",	-- Hex Addr	48C6	18630
x"00",	-- Hex Addr	48C7	18631
x"00",	-- Hex Addr	48C8	18632
x"00",	-- Hex Addr	48C9	18633
x"00",	-- Hex Addr	48CA	18634
x"00",	-- Hex Addr	48CB	18635
x"00",	-- Hex Addr	48CC	18636
x"00",	-- Hex Addr	48CD	18637
x"00",	-- Hex Addr	48CE	18638
x"00",	-- Hex Addr	48CF	18639
x"00",	-- Hex Addr	48D0	18640
x"00",	-- Hex Addr	48D1	18641
x"00",	-- Hex Addr	48D2	18642
x"00",	-- Hex Addr	48D3	18643
x"00",	-- Hex Addr	48D4	18644
x"00",	-- Hex Addr	48D5	18645
x"00",	-- Hex Addr	48D6	18646
x"00",	-- Hex Addr	48D7	18647
x"00",	-- Hex Addr	48D8	18648
x"00",	-- Hex Addr	48D9	18649
x"00",	-- Hex Addr	48DA	18650
x"00",	-- Hex Addr	48DB	18651
x"00",	-- Hex Addr	48DC	18652
x"00",	-- Hex Addr	48DD	18653
x"00",	-- Hex Addr	48DE	18654
x"00",	-- Hex Addr	48DF	18655
x"00",	-- Hex Addr	48E0	18656
x"00",	-- Hex Addr	48E1	18657
x"00",	-- Hex Addr	48E2	18658
x"00",	-- Hex Addr	48E3	18659
x"00",	-- Hex Addr	48E4	18660
x"00",	-- Hex Addr	48E5	18661
x"00",	-- Hex Addr	48E6	18662
x"00",	-- Hex Addr	48E7	18663
x"00",	-- Hex Addr	48E8	18664
x"00",	-- Hex Addr	48E9	18665
x"00",	-- Hex Addr	48EA	18666
x"00",	-- Hex Addr	48EB	18667
x"00",	-- Hex Addr	48EC	18668
x"00",	-- Hex Addr	48ED	18669
x"00",	-- Hex Addr	48EE	18670
x"00",	-- Hex Addr	48EF	18671
x"00",	-- Hex Addr	48F0	18672
x"00",	-- Hex Addr	48F1	18673
x"00",	-- Hex Addr	48F2	18674
x"00",	-- Hex Addr	48F3	18675
x"00",	-- Hex Addr	48F4	18676
x"00",	-- Hex Addr	48F5	18677
x"00",	-- Hex Addr	48F6	18678
x"00",	-- Hex Addr	48F7	18679
x"00",	-- Hex Addr	48F8	18680
x"00",	-- Hex Addr	48F9	18681
x"00",	-- Hex Addr	48FA	18682
x"00",	-- Hex Addr	48FB	18683
x"00",	-- Hex Addr	48FC	18684
x"00",	-- Hex Addr	48FD	18685
x"00",	-- Hex Addr	48FE	18686
x"00",	-- Hex Addr	48FF	18687
x"00",	-- Hex Addr	4900	18688
x"00",	-- Hex Addr	4901	18689
x"00",	-- Hex Addr	4902	18690
x"00",	-- Hex Addr	4903	18691
x"00",	-- Hex Addr	4904	18692
x"00",	-- Hex Addr	4905	18693
x"00",	-- Hex Addr	4906	18694
x"00",	-- Hex Addr	4907	18695
x"00",	-- Hex Addr	4908	18696
x"00",	-- Hex Addr	4909	18697
x"00",	-- Hex Addr	490A	18698
x"00",	-- Hex Addr	490B	18699
x"00",	-- Hex Addr	490C	18700
x"00",	-- Hex Addr	490D	18701
x"00",	-- Hex Addr	490E	18702
x"00",	-- Hex Addr	490F	18703
x"00",	-- Hex Addr	4910	18704
x"00",	-- Hex Addr	4911	18705
x"00",	-- Hex Addr	4912	18706
x"00",	-- Hex Addr	4913	18707
x"00",	-- Hex Addr	4914	18708
x"00",	-- Hex Addr	4915	18709
x"00",	-- Hex Addr	4916	18710
x"00",	-- Hex Addr	4917	18711
x"00",	-- Hex Addr	4918	18712
x"00",	-- Hex Addr	4919	18713
x"00",	-- Hex Addr	491A	18714
x"00",	-- Hex Addr	491B	18715
x"00",	-- Hex Addr	491C	18716
x"00",	-- Hex Addr	491D	18717
x"00",	-- Hex Addr	491E	18718
x"00",	-- Hex Addr	491F	18719
x"00",	-- Hex Addr	4920	18720
x"00",	-- Hex Addr	4921	18721
x"00",	-- Hex Addr	4922	18722
x"00",	-- Hex Addr	4923	18723
x"00",	-- Hex Addr	4924	18724
x"00",	-- Hex Addr	4925	18725
x"00",	-- Hex Addr	4926	18726
x"00",	-- Hex Addr	4927	18727
x"00",	-- Hex Addr	4928	18728
x"00",	-- Hex Addr	4929	18729
x"00",	-- Hex Addr	492A	18730
x"00",	-- Hex Addr	492B	18731
x"00",	-- Hex Addr	492C	18732
x"00",	-- Hex Addr	492D	18733
x"00",	-- Hex Addr	492E	18734
x"00",	-- Hex Addr	492F	18735
x"00",	-- Hex Addr	4930	18736
x"00",	-- Hex Addr	4931	18737
x"00",	-- Hex Addr	4932	18738
x"00",	-- Hex Addr	4933	18739
x"00",	-- Hex Addr	4934	18740
x"00",	-- Hex Addr	4935	18741
x"00",	-- Hex Addr	4936	18742
x"00",	-- Hex Addr	4937	18743
x"00",	-- Hex Addr	4938	18744
x"00",	-- Hex Addr	4939	18745
x"00",	-- Hex Addr	493A	18746
x"00",	-- Hex Addr	493B	18747
x"00",	-- Hex Addr	493C	18748
x"00",	-- Hex Addr	493D	18749
x"00",	-- Hex Addr	493E	18750
x"00",	-- Hex Addr	493F	18751
x"00",	-- Hex Addr	4940	18752
x"00",	-- Hex Addr	4941	18753
x"00",	-- Hex Addr	4942	18754
x"00",	-- Hex Addr	4943	18755
x"00",	-- Hex Addr	4944	18756
x"00",	-- Hex Addr	4945	18757
x"00",	-- Hex Addr	4946	18758
x"00",	-- Hex Addr	4947	18759
x"00",	-- Hex Addr	4948	18760
x"00",	-- Hex Addr	4949	18761
x"00",	-- Hex Addr	494A	18762
x"00",	-- Hex Addr	494B	18763
x"00",	-- Hex Addr	494C	18764
x"00",	-- Hex Addr	494D	18765
x"00",	-- Hex Addr	494E	18766
x"00",	-- Hex Addr	494F	18767
x"00",	-- Hex Addr	4950	18768
x"00",	-- Hex Addr	4951	18769
x"00",	-- Hex Addr	4952	18770
x"00",	-- Hex Addr	4953	18771
x"00",	-- Hex Addr	4954	18772
x"00",	-- Hex Addr	4955	18773
x"00",	-- Hex Addr	4956	18774
x"00",	-- Hex Addr	4957	18775
x"00",	-- Hex Addr	4958	18776
x"00",	-- Hex Addr	4959	18777
x"00",	-- Hex Addr	495A	18778
x"00",	-- Hex Addr	495B	18779
x"00",	-- Hex Addr	495C	18780
x"00",	-- Hex Addr	495D	18781
x"00",	-- Hex Addr	495E	18782
x"00",	-- Hex Addr	495F	18783
x"00",	-- Hex Addr	4960	18784
x"00",	-- Hex Addr	4961	18785
x"00",	-- Hex Addr	4962	18786
x"00",	-- Hex Addr	4963	18787
x"00",	-- Hex Addr	4964	18788
x"00",	-- Hex Addr	4965	18789
x"00",	-- Hex Addr	4966	18790
x"00",	-- Hex Addr	4967	18791
x"00",	-- Hex Addr	4968	18792
x"00",	-- Hex Addr	4969	18793
x"00",	-- Hex Addr	496A	18794
x"00",	-- Hex Addr	496B	18795
x"00",	-- Hex Addr	496C	18796
x"00",	-- Hex Addr	496D	18797
x"00",	-- Hex Addr	496E	18798
x"00",	-- Hex Addr	496F	18799
x"00",	-- Hex Addr	4970	18800
x"00",	-- Hex Addr	4971	18801
x"00",	-- Hex Addr	4972	18802
x"00",	-- Hex Addr	4973	18803
x"00",	-- Hex Addr	4974	18804
x"00",	-- Hex Addr	4975	18805
x"00",	-- Hex Addr	4976	18806
x"00",	-- Hex Addr	4977	18807
x"00",	-- Hex Addr	4978	18808
x"00",	-- Hex Addr	4979	18809
x"00",	-- Hex Addr	497A	18810
x"00",	-- Hex Addr	497B	18811
x"00",	-- Hex Addr	497C	18812
x"00",	-- Hex Addr	497D	18813
x"00",	-- Hex Addr	497E	18814
x"00",	-- Hex Addr	497F	18815
x"00",	-- Hex Addr	4980	18816
x"00",	-- Hex Addr	4981	18817
x"00",	-- Hex Addr	4982	18818
x"00",	-- Hex Addr	4983	18819
x"00",	-- Hex Addr	4984	18820
x"00",	-- Hex Addr	4985	18821
x"00",	-- Hex Addr	4986	18822
x"00",	-- Hex Addr	4987	18823
x"00",	-- Hex Addr	4988	18824
x"00",	-- Hex Addr	4989	18825
x"00",	-- Hex Addr	498A	18826
x"00",	-- Hex Addr	498B	18827
x"00",	-- Hex Addr	498C	18828
x"00",	-- Hex Addr	498D	18829
x"00",	-- Hex Addr	498E	18830
x"00",	-- Hex Addr	498F	18831
x"00",	-- Hex Addr	4990	18832
x"00",	-- Hex Addr	4991	18833
x"00",	-- Hex Addr	4992	18834
x"00",	-- Hex Addr	4993	18835
x"00",	-- Hex Addr	4994	18836
x"00",	-- Hex Addr	4995	18837
x"00",	-- Hex Addr	4996	18838
x"00",	-- Hex Addr	4997	18839
x"00",	-- Hex Addr	4998	18840
x"00",	-- Hex Addr	4999	18841
x"00",	-- Hex Addr	499A	18842
x"00",	-- Hex Addr	499B	18843
x"00",	-- Hex Addr	499C	18844
x"00",	-- Hex Addr	499D	18845
x"00",	-- Hex Addr	499E	18846
x"00",	-- Hex Addr	499F	18847
x"00",	-- Hex Addr	49A0	18848
x"00",	-- Hex Addr	49A1	18849
x"00",	-- Hex Addr	49A2	18850
x"00",	-- Hex Addr	49A3	18851
x"00",	-- Hex Addr	49A4	18852
x"00",	-- Hex Addr	49A5	18853
x"00",	-- Hex Addr	49A6	18854
x"00",	-- Hex Addr	49A7	18855
x"00",	-- Hex Addr	49A8	18856
x"00",	-- Hex Addr	49A9	18857
x"00",	-- Hex Addr	49AA	18858
x"00",	-- Hex Addr	49AB	18859
x"00",	-- Hex Addr	49AC	18860
x"00",	-- Hex Addr	49AD	18861
x"00",	-- Hex Addr	49AE	18862
x"00",	-- Hex Addr	49AF	18863
x"00",	-- Hex Addr	49B0	18864
x"00",	-- Hex Addr	49B1	18865
x"00",	-- Hex Addr	49B2	18866
x"00",	-- Hex Addr	49B3	18867
x"00",	-- Hex Addr	49B4	18868
x"00",	-- Hex Addr	49B5	18869
x"00",	-- Hex Addr	49B6	18870
x"00",	-- Hex Addr	49B7	18871
x"00",	-- Hex Addr	49B8	18872
x"00",	-- Hex Addr	49B9	18873
x"00",	-- Hex Addr	49BA	18874
x"00",	-- Hex Addr	49BB	18875
x"00",	-- Hex Addr	49BC	18876
x"00",	-- Hex Addr	49BD	18877
x"00",	-- Hex Addr	49BE	18878
x"00",	-- Hex Addr	49BF	18879
x"00",	-- Hex Addr	49C0	18880
x"00",	-- Hex Addr	49C1	18881
x"00",	-- Hex Addr	49C2	18882
x"00",	-- Hex Addr	49C3	18883
x"00",	-- Hex Addr	49C4	18884
x"00",	-- Hex Addr	49C5	18885
x"00",	-- Hex Addr	49C6	18886
x"00",	-- Hex Addr	49C7	18887
x"00",	-- Hex Addr	49C8	18888
x"00",	-- Hex Addr	49C9	18889
x"00",	-- Hex Addr	49CA	18890
x"00",	-- Hex Addr	49CB	18891
x"00",	-- Hex Addr	49CC	18892
x"00",	-- Hex Addr	49CD	18893
x"00",	-- Hex Addr	49CE	18894
x"00",	-- Hex Addr	49CF	18895
x"00",	-- Hex Addr	49D0	18896
x"00",	-- Hex Addr	49D1	18897
x"00",	-- Hex Addr	49D2	18898
x"00",	-- Hex Addr	49D3	18899
x"00",	-- Hex Addr	49D4	18900
x"00",	-- Hex Addr	49D5	18901
x"00",	-- Hex Addr	49D6	18902
x"00",	-- Hex Addr	49D7	18903
x"00",	-- Hex Addr	49D8	18904
x"00",	-- Hex Addr	49D9	18905
x"00",	-- Hex Addr	49DA	18906
x"00",	-- Hex Addr	49DB	18907
x"00",	-- Hex Addr	49DC	18908
x"00",	-- Hex Addr	49DD	18909
x"00",	-- Hex Addr	49DE	18910
x"00",	-- Hex Addr	49DF	18911
x"00",	-- Hex Addr	49E0	18912
x"00",	-- Hex Addr	49E1	18913
x"00",	-- Hex Addr	49E2	18914
x"00",	-- Hex Addr	49E3	18915
x"00",	-- Hex Addr	49E4	18916
x"00",	-- Hex Addr	49E5	18917
x"00",	-- Hex Addr	49E6	18918
x"00",	-- Hex Addr	49E7	18919
x"00",	-- Hex Addr	49E8	18920
x"00",	-- Hex Addr	49E9	18921
x"00",	-- Hex Addr	49EA	18922
x"00",	-- Hex Addr	49EB	18923
x"00",	-- Hex Addr	49EC	18924
x"00",	-- Hex Addr	49ED	18925
x"00",	-- Hex Addr	49EE	18926
x"00",	-- Hex Addr	49EF	18927
x"00",	-- Hex Addr	49F0	18928
x"00",	-- Hex Addr	49F1	18929
x"00",	-- Hex Addr	49F2	18930
x"00",	-- Hex Addr	49F3	18931
x"00",	-- Hex Addr	49F4	18932
x"00",	-- Hex Addr	49F5	18933
x"00",	-- Hex Addr	49F6	18934
x"00",	-- Hex Addr	49F7	18935
x"00",	-- Hex Addr	49F8	18936
x"00",	-- Hex Addr	49F9	18937
x"00",	-- Hex Addr	49FA	18938
x"00",	-- Hex Addr	49FB	18939
x"00",	-- Hex Addr	49FC	18940
x"00",	-- Hex Addr	49FD	18941
x"00",	-- Hex Addr	49FE	18942
x"00",	-- Hex Addr	49FF	18943
x"00",	-- Hex Addr	4A00	18944
x"00",	-- Hex Addr	4A01	18945
x"00",	-- Hex Addr	4A02	18946
x"00",	-- Hex Addr	4A03	18947
x"00",	-- Hex Addr	4A04	18948
x"00",	-- Hex Addr	4A05	18949
x"00",	-- Hex Addr	4A06	18950
x"00",	-- Hex Addr	4A07	18951
x"00",	-- Hex Addr	4A08	18952
x"00",	-- Hex Addr	4A09	18953
x"00",	-- Hex Addr	4A0A	18954
x"00",	-- Hex Addr	4A0B	18955
x"00",	-- Hex Addr	4A0C	18956
x"00",	-- Hex Addr	4A0D	18957
x"00",	-- Hex Addr	4A0E	18958
x"00",	-- Hex Addr	4A0F	18959
x"00",	-- Hex Addr	4A10	18960
x"00",	-- Hex Addr	4A11	18961
x"00",	-- Hex Addr	4A12	18962
x"00",	-- Hex Addr	4A13	18963
x"00",	-- Hex Addr	4A14	18964
x"00",	-- Hex Addr	4A15	18965
x"00",	-- Hex Addr	4A16	18966
x"00",	-- Hex Addr	4A17	18967
x"00",	-- Hex Addr	4A18	18968
x"00",	-- Hex Addr	4A19	18969
x"00",	-- Hex Addr	4A1A	18970
x"00",	-- Hex Addr	4A1B	18971
x"00",	-- Hex Addr	4A1C	18972
x"00",	-- Hex Addr	4A1D	18973
x"00",	-- Hex Addr	4A1E	18974
x"00",	-- Hex Addr	4A1F	18975
x"00",	-- Hex Addr	4A20	18976
x"00",	-- Hex Addr	4A21	18977
x"00",	-- Hex Addr	4A22	18978
x"00",	-- Hex Addr	4A23	18979
x"00",	-- Hex Addr	4A24	18980
x"00",	-- Hex Addr	4A25	18981
x"00",	-- Hex Addr	4A26	18982
x"00",	-- Hex Addr	4A27	18983
x"00",	-- Hex Addr	4A28	18984
x"00",	-- Hex Addr	4A29	18985
x"00",	-- Hex Addr	4A2A	18986
x"00",	-- Hex Addr	4A2B	18987
x"00",	-- Hex Addr	4A2C	18988
x"00",	-- Hex Addr	4A2D	18989
x"00",	-- Hex Addr	4A2E	18990
x"00",	-- Hex Addr	4A2F	18991
x"00",	-- Hex Addr	4A30	18992
x"00",	-- Hex Addr	4A31	18993
x"00",	-- Hex Addr	4A32	18994
x"00",	-- Hex Addr	4A33	18995
x"00",	-- Hex Addr	4A34	18996
x"00",	-- Hex Addr	4A35	18997
x"00",	-- Hex Addr	4A36	18998
x"00",	-- Hex Addr	4A37	18999
x"00",	-- Hex Addr	4A38	19000
x"00",	-- Hex Addr	4A39	19001
x"00",	-- Hex Addr	4A3A	19002
x"00",	-- Hex Addr	4A3B	19003
x"00",	-- Hex Addr	4A3C	19004
x"00",	-- Hex Addr	4A3D	19005
x"00",	-- Hex Addr	4A3E	19006
x"00",	-- Hex Addr	4A3F	19007
x"00",	-- Hex Addr	4A40	19008
x"00",	-- Hex Addr	4A41	19009
x"00",	-- Hex Addr	4A42	19010
x"00",	-- Hex Addr	4A43	19011
x"00",	-- Hex Addr	4A44	19012
x"00",	-- Hex Addr	4A45	19013
x"00",	-- Hex Addr	4A46	19014
x"00",	-- Hex Addr	4A47	19015
x"00",	-- Hex Addr	4A48	19016
x"00",	-- Hex Addr	4A49	19017
x"00",	-- Hex Addr	4A4A	19018
x"00",	-- Hex Addr	4A4B	19019
x"00",	-- Hex Addr	4A4C	19020
x"00",	-- Hex Addr	4A4D	19021
x"00",	-- Hex Addr	4A4E	19022
x"00",	-- Hex Addr	4A4F	19023
x"00",	-- Hex Addr	4A50	19024
x"00",	-- Hex Addr	4A51	19025
x"00",	-- Hex Addr	4A52	19026
x"00",	-- Hex Addr	4A53	19027
x"00",	-- Hex Addr	4A54	19028
x"00",	-- Hex Addr	4A55	19029
x"00",	-- Hex Addr	4A56	19030
x"00",	-- Hex Addr	4A57	19031
x"00",	-- Hex Addr	4A58	19032
x"00",	-- Hex Addr	4A59	19033
x"00",	-- Hex Addr	4A5A	19034
x"00",	-- Hex Addr	4A5B	19035
x"00",	-- Hex Addr	4A5C	19036
x"00",	-- Hex Addr	4A5D	19037
x"00",	-- Hex Addr	4A5E	19038
x"00",	-- Hex Addr	4A5F	19039
x"00",	-- Hex Addr	4A60	19040
x"00",	-- Hex Addr	4A61	19041
x"00",	-- Hex Addr	4A62	19042
x"00",	-- Hex Addr	4A63	19043
x"00",	-- Hex Addr	4A64	19044
x"00",	-- Hex Addr	4A65	19045
x"00",	-- Hex Addr	4A66	19046
x"00",	-- Hex Addr	4A67	19047
x"00",	-- Hex Addr	4A68	19048
x"00",	-- Hex Addr	4A69	19049
x"00",	-- Hex Addr	4A6A	19050
x"00",	-- Hex Addr	4A6B	19051
x"00",	-- Hex Addr	4A6C	19052
x"00",	-- Hex Addr	4A6D	19053
x"00",	-- Hex Addr	4A6E	19054
x"00",	-- Hex Addr	4A6F	19055
x"00",	-- Hex Addr	4A70	19056
x"00",	-- Hex Addr	4A71	19057
x"00",	-- Hex Addr	4A72	19058
x"00",	-- Hex Addr	4A73	19059
x"00",	-- Hex Addr	4A74	19060
x"00",	-- Hex Addr	4A75	19061
x"00",	-- Hex Addr	4A76	19062
x"00",	-- Hex Addr	4A77	19063
x"00",	-- Hex Addr	4A78	19064
x"00",	-- Hex Addr	4A79	19065
x"00",	-- Hex Addr	4A7A	19066
x"00",	-- Hex Addr	4A7B	19067
x"00",	-- Hex Addr	4A7C	19068
x"00",	-- Hex Addr	4A7D	19069
x"00",	-- Hex Addr	4A7E	19070
x"00",	-- Hex Addr	4A7F	19071
x"00",	-- Hex Addr	4A80	19072
x"00",	-- Hex Addr	4A81	19073
x"00",	-- Hex Addr	4A82	19074
x"00",	-- Hex Addr	4A83	19075
x"00",	-- Hex Addr	4A84	19076
x"00",	-- Hex Addr	4A85	19077
x"00",	-- Hex Addr	4A86	19078
x"00",	-- Hex Addr	4A87	19079
x"00",	-- Hex Addr	4A88	19080
x"00",	-- Hex Addr	4A89	19081
x"00",	-- Hex Addr	4A8A	19082
x"00",	-- Hex Addr	4A8B	19083
x"00",	-- Hex Addr	4A8C	19084
x"00",	-- Hex Addr	4A8D	19085
x"00",	-- Hex Addr	4A8E	19086
x"00",	-- Hex Addr	4A8F	19087
x"00",	-- Hex Addr	4A90	19088
x"00",	-- Hex Addr	4A91	19089
x"00",	-- Hex Addr	4A92	19090
x"00",	-- Hex Addr	4A93	19091
x"00",	-- Hex Addr	4A94	19092
x"00",	-- Hex Addr	4A95	19093
x"00",	-- Hex Addr	4A96	19094
x"00",	-- Hex Addr	4A97	19095
x"00",	-- Hex Addr	4A98	19096
x"00",	-- Hex Addr	4A99	19097
x"00",	-- Hex Addr	4A9A	19098
x"00",	-- Hex Addr	4A9B	19099
x"00",	-- Hex Addr	4A9C	19100
x"00",	-- Hex Addr	4A9D	19101
x"00",	-- Hex Addr	4A9E	19102
x"00",	-- Hex Addr	4A9F	19103
x"00",	-- Hex Addr	4AA0	19104
x"00",	-- Hex Addr	4AA1	19105
x"00",	-- Hex Addr	4AA2	19106
x"00",	-- Hex Addr	4AA3	19107
x"00",	-- Hex Addr	4AA4	19108
x"00",	-- Hex Addr	4AA5	19109
x"00",	-- Hex Addr	4AA6	19110
x"00",	-- Hex Addr	4AA7	19111
x"00",	-- Hex Addr	4AA8	19112
x"00",	-- Hex Addr	4AA9	19113
x"00",	-- Hex Addr	4AAA	19114
x"00",	-- Hex Addr	4AAB	19115
x"00",	-- Hex Addr	4AAC	19116
x"00",	-- Hex Addr	4AAD	19117
x"00",	-- Hex Addr	4AAE	19118
x"00",	-- Hex Addr	4AAF	19119
x"00",	-- Hex Addr	4AB0	19120
x"00",	-- Hex Addr	4AB1	19121
x"00",	-- Hex Addr	4AB2	19122
x"00",	-- Hex Addr	4AB3	19123
x"00",	-- Hex Addr	4AB4	19124
x"00",	-- Hex Addr	4AB5	19125
x"00",	-- Hex Addr	4AB6	19126
x"00",	-- Hex Addr	4AB7	19127
x"00",	-- Hex Addr	4AB8	19128
x"00",	-- Hex Addr	4AB9	19129
x"00",	-- Hex Addr	4ABA	19130
x"00",	-- Hex Addr	4ABB	19131
x"00",	-- Hex Addr	4ABC	19132
x"00",	-- Hex Addr	4ABD	19133
x"00",	-- Hex Addr	4ABE	19134
x"00",	-- Hex Addr	4ABF	19135
x"00",	-- Hex Addr	4AC0	19136
x"00",	-- Hex Addr	4AC1	19137
x"00",	-- Hex Addr	4AC2	19138
x"00",	-- Hex Addr	4AC3	19139
x"00",	-- Hex Addr	4AC4	19140
x"00",	-- Hex Addr	4AC5	19141
x"00",	-- Hex Addr	4AC6	19142
x"00",	-- Hex Addr	4AC7	19143
x"00",	-- Hex Addr	4AC8	19144
x"00",	-- Hex Addr	4AC9	19145
x"00",	-- Hex Addr	4ACA	19146
x"00",	-- Hex Addr	4ACB	19147
x"00",	-- Hex Addr	4ACC	19148
x"00",	-- Hex Addr	4ACD	19149
x"00",	-- Hex Addr	4ACE	19150
x"00",	-- Hex Addr	4ACF	19151
x"00",	-- Hex Addr	4AD0	19152
x"00",	-- Hex Addr	4AD1	19153
x"00",	-- Hex Addr	4AD2	19154
x"00",	-- Hex Addr	4AD3	19155
x"00",	-- Hex Addr	4AD4	19156
x"00",	-- Hex Addr	4AD5	19157
x"00",	-- Hex Addr	4AD6	19158
x"00",	-- Hex Addr	4AD7	19159
x"00",	-- Hex Addr	4AD8	19160
x"00",	-- Hex Addr	4AD9	19161
x"00",	-- Hex Addr	4ADA	19162
x"00",	-- Hex Addr	4ADB	19163
x"00",	-- Hex Addr	4ADC	19164
x"00",	-- Hex Addr	4ADD	19165
x"00",	-- Hex Addr	4ADE	19166
x"00",	-- Hex Addr	4ADF	19167
x"00",	-- Hex Addr	4AE0	19168
x"00",	-- Hex Addr	4AE1	19169
x"00",	-- Hex Addr	4AE2	19170
x"00",	-- Hex Addr	4AE3	19171
x"00",	-- Hex Addr	4AE4	19172
x"00",	-- Hex Addr	4AE5	19173
x"00",	-- Hex Addr	4AE6	19174
x"00",	-- Hex Addr	4AE7	19175
x"00",	-- Hex Addr	4AE8	19176
x"00",	-- Hex Addr	4AE9	19177
x"00",	-- Hex Addr	4AEA	19178
x"00",	-- Hex Addr	4AEB	19179
x"00",	-- Hex Addr	4AEC	19180
x"00",	-- Hex Addr	4AED	19181
x"00",	-- Hex Addr	4AEE	19182
x"00",	-- Hex Addr	4AEF	19183
x"00",	-- Hex Addr	4AF0	19184
x"00",	-- Hex Addr	4AF1	19185
x"00",	-- Hex Addr	4AF2	19186
x"00",	-- Hex Addr	4AF3	19187
x"00",	-- Hex Addr	4AF4	19188
x"00",	-- Hex Addr	4AF5	19189
x"00",	-- Hex Addr	4AF6	19190
x"00",	-- Hex Addr	4AF7	19191
x"00",	-- Hex Addr	4AF8	19192
x"00",	-- Hex Addr	4AF9	19193
x"00",	-- Hex Addr	4AFA	19194
x"00",	-- Hex Addr	4AFB	19195
x"00",	-- Hex Addr	4AFC	19196
x"00",	-- Hex Addr	4AFD	19197
x"00",	-- Hex Addr	4AFE	19198
x"00",	-- Hex Addr	4AFF	19199
x"00",	-- Hex Addr	4B00	19200
x"00",	-- Hex Addr	4B01	19201
x"00",	-- Hex Addr	4B02	19202
x"00",	-- Hex Addr	4B03	19203
x"00",	-- Hex Addr	4B04	19204
x"00",	-- Hex Addr	4B05	19205
x"00",	-- Hex Addr	4B06	19206
x"00",	-- Hex Addr	4B07	19207
x"00",	-- Hex Addr	4B08	19208
x"00",	-- Hex Addr	4B09	19209
x"00",	-- Hex Addr	4B0A	19210
x"00",	-- Hex Addr	4B0B	19211
x"00",	-- Hex Addr	4B0C	19212
x"00",	-- Hex Addr	4B0D	19213
x"00",	-- Hex Addr	4B0E	19214
x"00",	-- Hex Addr	4B0F	19215
x"00",	-- Hex Addr	4B10	19216
x"00",	-- Hex Addr	4B11	19217
x"00",	-- Hex Addr	4B12	19218
x"00",	-- Hex Addr	4B13	19219
x"00",	-- Hex Addr	4B14	19220
x"00",	-- Hex Addr	4B15	19221
x"00",	-- Hex Addr	4B16	19222
x"00",	-- Hex Addr	4B17	19223
x"00",	-- Hex Addr	4B18	19224
x"00",	-- Hex Addr	4B19	19225
x"00",	-- Hex Addr	4B1A	19226
x"00",	-- Hex Addr	4B1B	19227
x"00",	-- Hex Addr	4B1C	19228
x"00",	-- Hex Addr	4B1D	19229
x"00",	-- Hex Addr	4B1E	19230
x"00",	-- Hex Addr	4B1F	19231
x"00",	-- Hex Addr	4B20	19232
x"00",	-- Hex Addr	4B21	19233
x"00",	-- Hex Addr	4B22	19234
x"00",	-- Hex Addr	4B23	19235
x"00",	-- Hex Addr	4B24	19236
x"00",	-- Hex Addr	4B25	19237
x"00",	-- Hex Addr	4B26	19238
x"00",	-- Hex Addr	4B27	19239
x"00",	-- Hex Addr	4B28	19240
x"00",	-- Hex Addr	4B29	19241
x"00",	-- Hex Addr	4B2A	19242
x"00",	-- Hex Addr	4B2B	19243
x"00",	-- Hex Addr	4B2C	19244
x"00",	-- Hex Addr	4B2D	19245
x"00",	-- Hex Addr	4B2E	19246
x"00",	-- Hex Addr	4B2F	19247
x"00",	-- Hex Addr	4B30	19248
x"00",	-- Hex Addr	4B31	19249
x"00",	-- Hex Addr	4B32	19250
x"00",	-- Hex Addr	4B33	19251
x"00",	-- Hex Addr	4B34	19252
x"00",	-- Hex Addr	4B35	19253
x"00",	-- Hex Addr	4B36	19254
x"00",	-- Hex Addr	4B37	19255
x"00",	-- Hex Addr	4B38	19256
x"00",	-- Hex Addr	4B39	19257
x"00",	-- Hex Addr	4B3A	19258
x"00",	-- Hex Addr	4B3B	19259
x"00",	-- Hex Addr	4B3C	19260
x"00",	-- Hex Addr	4B3D	19261
x"00",	-- Hex Addr	4B3E	19262
x"00",	-- Hex Addr	4B3F	19263
x"00",	-- Hex Addr	4B40	19264
x"00",	-- Hex Addr	4B41	19265
x"00",	-- Hex Addr	4B42	19266
x"00",	-- Hex Addr	4B43	19267
x"00",	-- Hex Addr	4B44	19268
x"00",	-- Hex Addr	4B45	19269
x"00",	-- Hex Addr	4B46	19270
x"00",	-- Hex Addr	4B47	19271
x"00",	-- Hex Addr	4B48	19272
x"00",	-- Hex Addr	4B49	19273
x"00",	-- Hex Addr	4B4A	19274
x"00",	-- Hex Addr	4B4B	19275
x"00",	-- Hex Addr	4B4C	19276
x"00",	-- Hex Addr	4B4D	19277
x"00",	-- Hex Addr	4B4E	19278
x"00",	-- Hex Addr	4B4F	19279
x"00",	-- Hex Addr	4B50	19280
x"00",	-- Hex Addr	4B51	19281
x"00",	-- Hex Addr	4B52	19282
x"00",	-- Hex Addr	4B53	19283
x"00",	-- Hex Addr	4B54	19284
x"00",	-- Hex Addr	4B55	19285
x"00",	-- Hex Addr	4B56	19286
x"00",	-- Hex Addr	4B57	19287
x"00",	-- Hex Addr	4B58	19288
x"00",	-- Hex Addr	4B59	19289
x"00",	-- Hex Addr	4B5A	19290
x"00",	-- Hex Addr	4B5B	19291
x"00",	-- Hex Addr	4B5C	19292
x"00",	-- Hex Addr	4B5D	19293
x"00",	-- Hex Addr	4B5E	19294
x"00",	-- Hex Addr	4B5F	19295
x"00",	-- Hex Addr	4B60	19296
x"00",	-- Hex Addr	4B61	19297
x"00",	-- Hex Addr	4B62	19298
x"00",	-- Hex Addr	4B63	19299
x"00",	-- Hex Addr	4B64	19300
x"00",	-- Hex Addr	4B65	19301
x"00",	-- Hex Addr	4B66	19302
x"00",	-- Hex Addr	4B67	19303
x"00",	-- Hex Addr	4B68	19304
x"00",	-- Hex Addr	4B69	19305
x"00",	-- Hex Addr	4B6A	19306
x"00",	-- Hex Addr	4B6B	19307
x"00",	-- Hex Addr	4B6C	19308
x"00",	-- Hex Addr	4B6D	19309
x"00",	-- Hex Addr	4B6E	19310
x"00",	-- Hex Addr	4B6F	19311
x"00",	-- Hex Addr	4B70	19312
x"00",	-- Hex Addr	4B71	19313
x"00",	-- Hex Addr	4B72	19314
x"00",	-- Hex Addr	4B73	19315
x"00",	-- Hex Addr	4B74	19316
x"00",	-- Hex Addr	4B75	19317
x"00",	-- Hex Addr	4B76	19318
x"00",	-- Hex Addr	4B77	19319
x"00",	-- Hex Addr	4B78	19320
x"00",	-- Hex Addr	4B79	19321
x"00",	-- Hex Addr	4B7A	19322
x"00",	-- Hex Addr	4B7B	19323
x"00",	-- Hex Addr	4B7C	19324
x"00",	-- Hex Addr	4B7D	19325
x"00",	-- Hex Addr	4B7E	19326
x"00",	-- Hex Addr	4B7F	19327
x"00",	-- Hex Addr	4B80	19328
x"00",	-- Hex Addr	4B81	19329
x"00",	-- Hex Addr	4B82	19330
x"00",	-- Hex Addr	4B83	19331
x"00",	-- Hex Addr	4B84	19332
x"00",	-- Hex Addr	4B85	19333
x"00",	-- Hex Addr	4B86	19334
x"00",	-- Hex Addr	4B87	19335
x"00",	-- Hex Addr	4B88	19336
x"00",	-- Hex Addr	4B89	19337
x"00",	-- Hex Addr	4B8A	19338
x"00",	-- Hex Addr	4B8B	19339
x"00",	-- Hex Addr	4B8C	19340
x"00",	-- Hex Addr	4B8D	19341
x"00",	-- Hex Addr	4B8E	19342
x"00",	-- Hex Addr	4B8F	19343
x"00",	-- Hex Addr	4B90	19344
x"00",	-- Hex Addr	4B91	19345
x"00",	-- Hex Addr	4B92	19346
x"00",	-- Hex Addr	4B93	19347
x"00",	-- Hex Addr	4B94	19348
x"00",	-- Hex Addr	4B95	19349
x"00",	-- Hex Addr	4B96	19350
x"00",	-- Hex Addr	4B97	19351
x"00",	-- Hex Addr	4B98	19352
x"00",	-- Hex Addr	4B99	19353
x"00",	-- Hex Addr	4B9A	19354
x"00",	-- Hex Addr	4B9B	19355
x"00",	-- Hex Addr	4B9C	19356
x"00",	-- Hex Addr	4B9D	19357
x"00",	-- Hex Addr	4B9E	19358
x"00",	-- Hex Addr	4B9F	19359
x"00",	-- Hex Addr	4BA0	19360
x"00",	-- Hex Addr	4BA1	19361
x"00",	-- Hex Addr	4BA2	19362
x"00",	-- Hex Addr	4BA3	19363
x"00",	-- Hex Addr	4BA4	19364
x"00",	-- Hex Addr	4BA5	19365
x"00",	-- Hex Addr	4BA6	19366
x"00",	-- Hex Addr	4BA7	19367
x"00",	-- Hex Addr	4BA8	19368
x"00",	-- Hex Addr	4BA9	19369
x"00",	-- Hex Addr	4BAA	19370
x"00",	-- Hex Addr	4BAB	19371
x"00",	-- Hex Addr	4BAC	19372
x"00",	-- Hex Addr	4BAD	19373
x"00",	-- Hex Addr	4BAE	19374
x"00",	-- Hex Addr	4BAF	19375
x"00",	-- Hex Addr	4BB0	19376
x"00",	-- Hex Addr	4BB1	19377
x"00",	-- Hex Addr	4BB2	19378
x"00",	-- Hex Addr	4BB3	19379
x"00",	-- Hex Addr	4BB4	19380
x"00",	-- Hex Addr	4BB5	19381
x"00",	-- Hex Addr	4BB6	19382
x"00",	-- Hex Addr	4BB7	19383
x"00",	-- Hex Addr	4BB8	19384
x"00",	-- Hex Addr	4BB9	19385
x"00",	-- Hex Addr	4BBA	19386
x"00",	-- Hex Addr	4BBB	19387
x"00",	-- Hex Addr	4BBC	19388
x"00",	-- Hex Addr	4BBD	19389
x"00",	-- Hex Addr	4BBE	19390
x"00",	-- Hex Addr	4BBF	19391
x"00",	-- Hex Addr	4BC0	19392
x"00",	-- Hex Addr	4BC1	19393
x"00",	-- Hex Addr	4BC2	19394
x"00",	-- Hex Addr	4BC3	19395
x"00",	-- Hex Addr	4BC4	19396
x"00",	-- Hex Addr	4BC5	19397
x"00",	-- Hex Addr	4BC6	19398
x"00",	-- Hex Addr	4BC7	19399
x"00",	-- Hex Addr	4BC8	19400
x"00",	-- Hex Addr	4BC9	19401
x"00",	-- Hex Addr	4BCA	19402
x"00",	-- Hex Addr	4BCB	19403
x"00",	-- Hex Addr	4BCC	19404
x"00",	-- Hex Addr	4BCD	19405
x"00",	-- Hex Addr	4BCE	19406
x"00",	-- Hex Addr	4BCF	19407
x"00",	-- Hex Addr	4BD0	19408
x"00",	-- Hex Addr	4BD1	19409
x"00",	-- Hex Addr	4BD2	19410
x"00",	-- Hex Addr	4BD3	19411
x"00",	-- Hex Addr	4BD4	19412
x"00",	-- Hex Addr	4BD5	19413
x"00",	-- Hex Addr	4BD6	19414
x"00",	-- Hex Addr	4BD7	19415
x"00",	-- Hex Addr	4BD8	19416
x"00",	-- Hex Addr	4BD9	19417
x"00",	-- Hex Addr	4BDA	19418
x"00",	-- Hex Addr	4BDB	19419
x"00",	-- Hex Addr	4BDC	19420
x"00",	-- Hex Addr	4BDD	19421
x"00",	-- Hex Addr	4BDE	19422
x"00",	-- Hex Addr	4BDF	19423
x"00",	-- Hex Addr	4BE0	19424
x"00",	-- Hex Addr	4BE1	19425
x"00",	-- Hex Addr	4BE2	19426
x"00",	-- Hex Addr	4BE3	19427
x"00",	-- Hex Addr	4BE4	19428
x"00",	-- Hex Addr	4BE5	19429
x"00",	-- Hex Addr	4BE6	19430
x"00",	-- Hex Addr	4BE7	19431
x"00",	-- Hex Addr	4BE8	19432
x"00",	-- Hex Addr	4BE9	19433
x"00",	-- Hex Addr	4BEA	19434
x"00",	-- Hex Addr	4BEB	19435
x"00",	-- Hex Addr	4BEC	19436
x"00",	-- Hex Addr	4BED	19437
x"00",	-- Hex Addr	4BEE	19438
x"00",	-- Hex Addr	4BEF	19439
x"00",	-- Hex Addr	4BF0	19440
x"00",	-- Hex Addr	4BF1	19441
x"00",	-- Hex Addr	4BF2	19442
x"00",	-- Hex Addr	4BF3	19443
x"00",	-- Hex Addr	4BF4	19444
x"00",	-- Hex Addr	4BF5	19445
x"00",	-- Hex Addr	4BF6	19446
x"00",	-- Hex Addr	4BF7	19447
x"00",	-- Hex Addr	4BF8	19448
x"00",	-- Hex Addr	4BF9	19449
x"00",	-- Hex Addr	4BFA	19450
x"00",	-- Hex Addr	4BFB	19451
x"00",	-- Hex Addr	4BFC	19452
x"00",	-- Hex Addr	4BFD	19453
x"00",	-- Hex Addr	4BFE	19454
x"00",	-- Hex Addr	4BFF	19455
x"00",	-- Hex Addr	4C00	19456
x"00",	-- Hex Addr	4C01	19457
x"00",	-- Hex Addr	4C02	19458
x"00",	-- Hex Addr	4C03	19459
x"00",	-- Hex Addr	4C04	19460
x"00",	-- Hex Addr	4C05	19461
x"00",	-- Hex Addr	4C06	19462
x"00",	-- Hex Addr	4C07	19463
x"00",	-- Hex Addr	4C08	19464
x"00",	-- Hex Addr	4C09	19465
x"00",	-- Hex Addr	4C0A	19466
x"00",	-- Hex Addr	4C0B	19467
x"00",	-- Hex Addr	4C0C	19468
x"00",	-- Hex Addr	4C0D	19469
x"00",	-- Hex Addr	4C0E	19470
x"00",	-- Hex Addr	4C0F	19471
x"00",	-- Hex Addr	4C10	19472
x"00",	-- Hex Addr	4C11	19473
x"00",	-- Hex Addr	4C12	19474
x"00",	-- Hex Addr	4C13	19475
x"00",	-- Hex Addr	4C14	19476
x"00",	-- Hex Addr	4C15	19477
x"00",	-- Hex Addr	4C16	19478
x"00",	-- Hex Addr	4C17	19479
x"00",	-- Hex Addr	4C18	19480
x"00",	-- Hex Addr	4C19	19481
x"00",	-- Hex Addr	4C1A	19482
x"00",	-- Hex Addr	4C1B	19483
x"00",	-- Hex Addr	4C1C	19484
x"00",	-- Hex Addr	4C1D	19485
x"00",	-- Hex Addr	4C1E	19486
x"00",	-- Hex Addr	4C1F	19487
x"00",	-- Hex Addr	4C20	19488
x"00",	-- Hex Addr	4C21	19489
x"00",	-- Hex Addr	4C22	19490
x"00",	-- Hex Addr	4C23	19491
x"00",	-- Hex Addr	4C24	19492
x"00",	-- Hex Addr	4C25	19493
x"00",	-- Hex Addr	4C26	19494
x"00",	-- Hex Addr	4C27	19495
x"00",	-- Hex Addr	4C28	19496
x"00",	-- Hex Addr	4C29	19497
x"00",	-- Hex Addr	4C2A	19498
x"00",	-- Hex Addr	4C2B	19499
x"00",	-- Hex Addr	4C2C	19500
x"00",	-- Hex Addr	4C2D	19501
x"00",	-- Hex Addr	4C2E	19502
x"00",	-- Hex Addr	4C2F	19503
x"00",	-- Hex Addr	4C30	19504
x"00",	-- Hex Addr	4C31	19505
x"00",	-- Hex Addr	4C32	19506
x"00",	-- Hex Addr	4C33	19507
x"00",	-- Hex Addr	4C34	19508
x"00",	-- Hex Addr	4C35	19509
x"00",	-- Hex Addr	4C36	19510
x"00",	-- Hex Addr	4C37	19511
x"00",	-- Hex Addr	4C38	19512
x"00",	-- Hex Addr	4C39	19513
x"00",	-- Hex Addr	4C3A	19514
x"00",	-- Hex Addr	4C3B	19515
x"00",	-- Hex Addr	4C3C	19516
x"00",	-- Hex Addr	4C3D	19517
x"00",	-- Hex Addr	4C3E	19518
x"00",	-- Hex Addr	4C3F	19519
x"00",	-- Hex Addr	4C40	19520
x"00",	-- Hex Addr	4C41	19521
x"00",	-- Hex Addr	4C42	19522
x"00",	-- Hex Addr	4C43	19523
x"00",	-- Hex Addr	4C44	19524
x"00",	-- Hex Addr	4C45	19525
x"00",	-- Hex Addr	4C46	19526
x"00",	-- Hex Addr	4C47	19527
x"00",	-- Hex Addr	4C48	19528
x"00",	-- Hex Addr	4C49	19529
x"00",	-- Hex Addr	4C4A	19530
x"00",	-- Hex Addr	4C4B	19531
x"00",	-- Hex Addr	4C4C	19532
x"00",	-- Hex Addr	4C4D	19533
x"00",	-- Hex Addr	4C4E	19534
x"00",	-- Hex Addr	4C4F	19535
x"00",	-- Hex Addr	4C50	19536
x"00",	-- Hex Addr	4C51	19537
x"00",	-- Hex Addr	4C52	19538
x"00",	-- Hex Addr	4C53	19539
x"00",	-- Hex Addr	4C54	19540
x"00",	-- Hex Addr	4C55	19541
x"00",	-- Hex Addr	4C56	19542
x"00",	-- Hex Addr	4C57	19543
x"00",	-- Hex Addr	4C58	19544
x"00",	-- Hex Addr	4C59	19545
x"00",	-- Hex Addr	4C5A	19546
x"00",	-- Hex Addr	4C5B	19547
x"00",	-- Hex Addr	4C5C	19548
x"00",	-- Hex Addr	4C5D	19549
x"00",	-- Hex Addr	4C5E	19550
x"00",	-- Hex Addr	4C5F	19551
x"00",	-- Hex Addr	4C60	19552
x"00",	-- Hex Addr	4C61	19553
x"00",	-- Hex Addr	4C62	19554
x"00",	-- Hex Addr	4C63	19555
x"00",	-- Hex Addr	4C64	19556
x"00",	-- Hex Addr	4C65	19557
x"00",	-- Hex Addr	4C66	19558
x"00",	-- Hex Addr	4C67	19559
x"00",	-- Hex Addr	4C68	19560
x"00",	-- Hex Addr	4C69	19561
x"00",	-- Hex Addr	4C6A	19562
x"00",	-- Hex Addr	4C6B	19563
x"00",	-- Hex Addr	4C6C	19564
x"00",	-- Hex Addr	4C6D	19565
x"00",	-- Hex Addr	4C6E	19566
x"00",	-- Hex Addr	4C6F	19567
x"00",	-- Hex Addr	4C70	19568
x"00",	-- Hex Addr	4C71	19569
x"00",	-- Hex Addr	4C72	19570
x"00",	-- Hex Addr	4C73	19571
x"00",	-- Hex Addr	4C74	19572
x"00",	-- Hex Addr	4C75	19573
x"00",	-- Hex Addr	4C76	19574
x"00",	-- Hex Addr	4C77	19575
x"00",	-- Hex Addr	4C78	19576
x"00",	-- Hex Addr	4C79	19577
x"00",	-- Hex Addr	4C7A	19578
x"00",	-- Hex Addr	4C7B	19579
x"00",	-- Hex Addr	4C7C	19580
x"00",	-- Hex Addr	4C7D	19581
x"00",	-- Hex Addr	4C7E	19582
x"00",	-- Hex Addr	4C7F	19583
x"00",	-- Hex Addr	4C80	19584
x"00",	-- Hex Addr	4C81	19585
x"00",	-- Hex Addr	4C82	19586
x"00",	-- Hex Addr	4C83	19587
x"00",	-- Hex Addr	4C84	19588
x"00",	-- Hex Addr	4C85	19589
x"00",	-- Hex Addr	4C86	19590
x"00",	-- Hex Addr	4C87	19591
x"00",	-- Hex Addr	4C88	19592
x"00",	-- Hex Addr	4C89	19593
x"00",	-- Hex Addr	4C8A	19594
x"00",	-- Hex Addr	4C8B	19595
x"00",	-- Hex Addr	4C8C	19596
x"00",	-- Hex Addr	4C8D	19597
x"00",	-- Hex Addr	4C8E	19598
x"00",	-- Hex Addr	4C8F	19599
x"00",	-- Hex Addr	4C90	19600
x"00",	-- Hex Addr	4C91	19601
x"00",	-- Hex Addr	4C92	19602
x"00",	-- Hex Addr	4C93	19603
x"00",	-- Hex Addr	4C94	19604
x"00",	-- Hex Addr	4C95	19605
x"00",	-- Hex Addr	4C96	19606
x"00",	-- Hex Addr	4C97	19607
x"00",	-- Hex Addr	4C98	19608
x"00",	-- Hex Addr	4C99	19609
x"00",	-- Hex Addr	4C9A	19610
x"00",	-- Hex Addr	4C9B	19611
x"00",	-- Hex Addr	4C9C	19612
x"00",	-- Hex Addr	4C9D	19613
x"00",	-- Hex Addr	4C9E	19614
x"00",	-- Hex Addr	4C9F	19615
x"00",	-- Hex Addr	4CA0	19616
x"00",	-- Hex Addr	4CA1	19617
x"00",	-- Hex Addr	4CA2	19618
x"00",	-- Hex Addr	4CA3	19619
x"00",	-- Hex Addr	4CA4	19620
x"00",	-- Hex Addr	4CA5	19621
x"00",	-- Hex Addr	4CA6	19622
x"00",	-- Hex Addr	4CA7	19623
x"00",	-- Hex Addr	4CA8	19624
x"00",	-- Hex Addr	4CA9	19625
x"00",	-- Hex Addr	4CAA	19626
x"00",	-- Hex Addr	4CAB	19627
x"00",	-- Hex Addr	4CAC	19628
x"00",	-- Hex Addr	4CAD	19629
x"00",	-- Hex Addr	4CAE	19630
x"00",	-- Hex Addr	4CAF	19631
x"00",	-- Hex Addr	4CB0	19632
x"00",	-- Hex Addr	4CB1	19633
x"00",	-- Hex Addr	4CB2	19634
x"00",	-- Hex Addr	4CB3	19635
x"00",	-- Hex Addr	4CB4	19636
x"00",	-- Hex Addr	4CB5	19637
x"00",	-- Hex Addr	4CB6	19638
x"00",	-- Hex Addr	4CB7	19639
x"00",	-- Hex Addr	4CB8	19640
x"00",	-- Hex Addr	4CB9	19641
x"00",	-- Hex Addr	4CBA	19642
x"00",	-- Hex Addr	4CBB	19643
x"00",	-- Hex Addr	4CBC	19644
x"00",	-- Hex Addr	4CBD	19645
x"00",	-- Hex Addr	4CBE	19646
x"00",	-- Hex Addr	4CBF	19647
x"00",	-- Hex Addr	4CC0	19648
x"00",	-- Hex Addr	4CC1	19649
x"00",	-- Hex Addr	4CC2	19650
x"00",	-- Hex Addr	4CC3	19651
x"00",	-- Hex Addr	4CC4	19652
x"00",	-- Hex Addr	4CC5	19653
x"00",	-- Hex Addr	4CC6	19654
x"00",	-- Hex Addr	4CC7	19655
x"00",	-- Hex Addr	4CC8	19656
x"00",	-- Hex Addr	4CC9	19657
x"00",	-- Hex Addr	4CCA	19658
x"00",	-- Hex Addr	4CCB	19659
x"00",	-- Hex Addr	4CCC	19660
x"00",	-- Hex Addr	4CCD	19661
x"00",	-- Hex Addr	4CCE	19662
x"00",	-- Hex Addr	4CCF	19663
x"00",	-- Hex Addr	4CD0	19664
x"00",	-- Hex Addr	4CD1	19665
x"00",	-- Hex Addr	4CD2	19666
x"00",	-- Hex Addr	4CD3	19667
x"00",	-- Hex Addr	4CD4	19668
x"00",	-- Hex Addr	4CD5	19669
x"00",	-- Hex Addr	4CD6	19670
x"00",	-- Hex Addr	4CD7	19671
x"00",	-- Hex Addr	4CD8	19672
x"00",	-- Hex Addr	4CD9	19673
x"00",	-- Hex Addr	4CDA	19674
x"00",	-- Hex Addr	4CDB	19675
x"00",	-- Hex Addr	4CDC	19676
x"00",	-- Hex Addr	4CDD	19677
x"00",	-- Hex Addr	4CDE	19678
x"00",	-- Hex Addr	4CDF	19679
x"00",	-- Hex Addr	4CE0	19680
x"00",	-- Hex Addr	4CE1	19681
x"00",	-- Hex Addr	4CE2	19682
x"00",	-- Hex Addr	4CE3	19683
x"00",	-- Hex Addr	4CE4	19684
x"00",	-- Hex Addr	4CE5	19685
x"00",	-- Hex Addr	4CE6	19686
x"00",	-- Hex Addr	4CE7	19687
x"00",	-- Hex Addr	4CE8	19688
x"00",	-- Hex Addr	4CE9	19689
x"00",	-- Hex Addr	4CEA	19690
x"00",	-- Hex Addr	4CEB	19691
x"00",	-- Hex Addr	4CEC	19692
x"00",	-- Hex Addr	4CED	19693
x"00",	-- Hex Addr	4CEE	19694
x"00",	-- Hex Addr	4CEF	19695
x"00",	-- Hex Addr	4CF0	19696
x"00",	-- Hex Addr	4CF1	19697
x"00",	-- Hex Addr	4CF2	19698
x"00",	-- Hex Addr	4CF3	19699
x"00",	-- Hex Addr	4CF4	19700
x"00",	-- Hex Addr	4CF5	19701
x"00",	-- Hex Addr	4CF6	19702
x"00",	-- Hex Addr	4CF7	19703
x"00",	-- Hex Addr	4CF8	19704
x"00",	-- Hex Addr	4CF9	19705
x"00",	-- Hex Addr	4CFA	19706
x"00",	-- Hex Addr	4CFB	19707
x"00",	-- Hex Addr	4CFC	19708
x"00",	-- Hex Addr	4CFD	19709
x"00",	-- Hex Addr	4CFE	19710
x"00",	-- Hex Addr	4CFF	19711
x"00",	-- Hex Addr	4D00	19712
x"00",	-- Hex Addr	4D01	19713
x"00",	-- Hex Addr	4D02	19714
x"00",	-- Hex Addr	4D03	19715
x"00",	-- Hex Addr	4D04	19716
x"00",	-- Hex Addr	4D05	19717
x"00",	-- Hex Addr	4D06	19718
x"00",	-- Hex Addr	4D07	19719
x"00",	-- Hex Addr	4D08	19720
x"00",	-- Hex Addr	4D09	19721
x"00",	-- Hex Addr	4D0A	19722
x"00",	-- Hex Addr	4D0B	19723
x"00",	-- Hex Addr	4D0C	19724
x"00",	-- Hex Addr	4D0D	19725
x"00",	-- Hex Addr	4D0E	19726
x"00",	-- Hex Addr	4D0F	19727
x"00",	-- Hex Addr	4D10	19728
x"00",	-- Hex Addr	4D11	19729
x"00",	-- Hex Addr	4D12	19730
x"00",	-- Hex Addr	4D13	19731
x"00",	-- Hex Addr	4D14	19732
x"00",	-- Hex Addr	4D15	19733
x"00",	-- Hex Addr	4D16	19734
x"00",	-- Hex Addr	4D17	19735
x"00",	-- Hex Addr	4D18	19736
x"00",	-- Hex Addr	4D19	19737
x"00",	-- Hex Addr	4D1A	19738
x"00",	-- Hex Addr	4D1B	19739
x"00",	-- Hex Addr	4D1C	19740
x"00",	-- Hex Addr	4D1D	19741
x"00",	-- Hex Addr	4D1E	19742
x"00",	-- Hex Addr	4D1F	19743
x"00",	-- Hex Addr	4D20	19744
x"00",	-- Hex Addr	4D21	19745
x"00",	-- Hex Addr	4D22	19746
x"00",	-- Hex Addr	4D23	19747
x"00",	-- Hex Addr	4D24	19748
x"00",	-- Hex Addr	4D25	19749
x"00",	-- Hex Addr	4D26	19750
x"00",	-- Hex Addr	4D27	19751
x"00",	-- Hex Addr	4D28	19752
x"00",	-- Hex Addr	4D29	19753
x"00",	-- Hex Addr	4D2A	19754
x"00",	-- Hex Addr	4D2B	19755
x"00",	-- Hex Addr	4D2C	19756
x"00",	-- Hex Addr	4D2D	19757
x"00",	-- Hex Addr	4D2E	19758
x"00",	-- Hex Addr	4D2F	19759
x"00",	-- Hex Addr	4D30	19760
x"00",	-- Hex Addr	4D31	19761
x"00",	-- Hex Addr	4D32	19762
x"00",	-- Hex Addr	4D33	19763
x"00",	-- Hex Addr	4D34	19764
x"00",	-- Hex Addr	4D35	19765
x"00",	-- Hex Addr	4D36	19766
x"00",	-- Hex Addr	4D37	19767
x"00",	-- Hex Addr	4D38	19768
x"00",	-- Hex Addr	4D39	19769
x"00",	-- Hex Addr	4D3A	19770
x"00",	-- Hex Addr	4D3B	19771
x"00",	-- Hex Addr	4D3C	19772
x"00",	-- Hex Addr	4D3D	19773
x"00",	-- Hex Addr	4D3E	19774
x"00",	-- Hex Addr	4D3F	19775
x"00",	-- Hex Addr	4D40	19776
x"00",	-- Hex Addr	4D41	19777
x"00",	-- Hex Addr	4D42	19778
x"00",	-- Hex Addr	4D43	19779
x"00",	-- Hex Addr	4D44	19780
x"00",	-- Hex Addr	4D45	19781
x"00",	-- Hex Addr	4D46	19782
x"00",	-- Hex Addr	4D47	19783
x"00",	-- Hex Addr	4D48	19784
x"00",	-- Hex Addr	4D49	19785
x"00",	-- Hex Addr	4D4A	19786
x"00",	-- Hex Addr	4D4B	19787
x"00",	-- Hex Addr	4D4C	19788
x"00",	-- Hex Addr	4D4D	19789
x"00",	-- Hex Addr	4D4E	19790
x"00",	-- Hex Addr	4D4F	19791
x"00",	-- Hex Addr	4D50	19792
x"00",	-- Hex Addr	4D51	19793
x"00",	-- Hex Addr	4D52	19794
x"00",	-- Hex Addr	4D53	19795
x"00",	-- Hex Addr	4D54	19796
x"00",	-- Hex Addr	4D55	19797
x"00",	-- Hex Addr	4D56	19798
x"00",	-- Hex Addr	4D57	19799
x"00",	-- Hex Addr	4D58	19800
x"00",	-- Hex Addr	4D59	19801
x"00",	-- Hex Addr	4D5A	19802
x"00",	-- Hex Addr	4D5B	19803
x"00",	-- Hex Addr	4D5C	19804
x"00",	-- Hex Addr	4D5D	19805
x"00",	-- Hex Addr	4D5E	19806
x"00",	-- Hex Addr	4D5F	19807
x"00",	-- Hex Addr	4D60	19808
x"00",	-- Hex Addr	4D61	19809
x"00",	-- Hex Addr	4D62	19810
x"00",	-- Hex Addr	4D63	19811
x"00",	-- Hex Addr	4D64	19812
x"00",	-- Hex Addr	4D65	19813
x"00",	-- Hex Addr	4D66	19814
x"00",	-- Hex Addr	4D67	19815
x"00",	-- Hex Addr	4D68	19816
x"00",	-- Hex Addr	4D69	19817
x"00",	-- Hex Addr	4D6A	19818
x"00",	-- Hex Addr	4D6B	19819
x"00",	-- Hex Addr	4D6C	19820
x"00",	-- Hex Addr	4D6D	19821
x"00",	-- Hex Addr	4D6E	19822
x"00",	-- Hex Addr	4D6F	19823
x"00",	-- Hex Addr	4D70	19824
x"00",	-- Hex Addr	4D71	19825
x"00",	-- Hex Addr	4D72	19826
x"00",	-- Hex Addr	4D73	19827
x"00",	-- Hex Addr	4D74	19828
x"00",	-- Hex Addr	4D75	19829
x"00",	-- Hex Addr	4D76	19830
x"00",	-- Hex Addr	4D77	19831
x"00",	-- Hex Addr	4D78	19832
x"00",	-- Hex Addr	4D79	19833
x"00",	-- Hex Addr	4D7A	19834
x"00",	-- Hex Addr	4D7B	19835
x"00",	-- Hex Addr	4D7C	19836
x"00",	-- Hex Addr	4D7D	19837
x"00",	-- Hex Addr	4D7E	19838
x"00",	-- Hex Addr	4D7F	19839
x"00",	-- Hex Addr	4D80	19840
x"00",	-- Hex Addr	4D81	19841
x"00",	-- Hex Addr	4D82	19842
x"00",	-- Hex Addr	4D83	19843
x"00",	-- Hex Addr	4D84	19844
x"00",	-- Hex Addr	4D85	19845
x"00",	-- Hex Addr	4D86	19846
x"00",	-- Hex Addr	4D87	19847
x"00",	-- Hex Addr	4D88	19848
x"00",	-- Hex Addr	4D89	19849
x"00",	-- Hex Addr	4D8A	19850
x"00",	-- Hex Addr	4D8B	19851
x"00",	-- Hex Addr	4D8C	19852
x"00",	-- Hex Addr	4D8D	19853
x"00",	-- Hex Addr	4D8E	19854
x"00",	-- Hex Addr	4D8F	19855
x"00",	-- Hex Addr	4D90	19856
x"00",	-- Hex Addr	4D91	19857
x"00",	-- Hex Addr	4D92	19858
x"00",	-- Hex Addr	4D93	19859
x"00",	-- Hex Addr	4D94	19860
x"00",	-- Hex Addr	4D95	19861
x"00",	-- Hex Addr	4D96	19862
x"00",	-- Hex Addr	4D97	19863
x"00",	-- Hex Addr	4D98	19864
x"00",	-- Hex Addr	4D99	19865
x"00",	-- Hex Addr	4D9A	19866
x"00",	-- Hex Addr	4D9B	19867
x"00",	-- Hex Addr	4D9C	19868
x"00",	-- Hex Addr	4D9D	19869
x"00",	-- Hex Addr	4D9E	19870
x"00",	-- Hex Addr	4D9F	19871
x"00",	-- Hex Addr	4DA0	19872
x"00",	-- Hex Addr	4DA1	19873
x"00",	-- Hex Addr	4DA2	19874
x"00",	-- Hex Addr	4DA3	19875
x"00",	-- Hex Addr	4DA4	19876
x"00",	-- Hex Addr	4DA5	19877
x"00",	-- Hex Addr	4DA6	19878
x"00",	-- Hex Addr	4DA7	19879
x"00",	-- Hex Addr	4DA8	19880
x"00",	-- Hex Addr	4DA9	19881
x"00",	-- Hex Addr	4DAA	19882
x"00",	-- Hex Addr	4DAB	19883
x"00",	-- Hex Addr	4DAC	19884
x"00",	-- Hex Addr	4DAD	19885
x"00",	-- Hex Addr	4DAE	19886
x"00",	-- Hex Addr	4DAF	19887
x"00",	-- Hex Addr	4DB0	19888
x"00",	-- Hex Addr	4DB1	19889
x"00",	-- Hex Addr	4DB2	19890
x"00",	-- Hex Addr	4DB3	19891
x"00",	-- Hex Addr	4DB4	19892
x"00",	-- Hex Addr	4DB5	19893
x"00",	-- Hex Addr	4DB6	19894
x"00",	-- Hex Addr	4DB7	19895
x"00",	-- Hex Addr	4DB8	19896
x"00",	-- Hex Addr	4DB9	19897
x"00",	-- Hex Addr	4DBA	19898
x"00",	-- Hex Addr	4DBB	19899
x"00",	-- Hex Addr	4DBC	19900
x"00",	-- Hex Addr	4DBD	19901
x"00",	-- Hex Addr	4DBE	19902
x"00",	-- Hex Addr	4DBF	19903
x"00",	-- Hex Addr	4DC0	19904
x"00",	-- Hex Addr	4DC1	19905
x"00",	-- Hex Addr	4DC2	19906
x"00",	-- Hex Addr	4DC3	19907
x"00",	-- Hex Addr	4DC4	19908
x"00",	-- Hex Addr	4DC5	19909
x"00",	-- Hex Addr	4DC6	19910
x"00",	-- Hex Addr	4DC7	19911
x"00",	-- Hex Addr	4DC8	19912
x"00",	-- Hex Addr	4DC9	19913
x"00",	-- Hex Addr	4DCA	19914
x"00",	-- Hex Addr	4DCB	19915
x"00",	-- Hex Addr	4DCC	19916
x"00",	-- Hex Addr	4DCD	19917
x"00",	-- Hex Addr	4DCE	19918
x"00",	-- Hex Addr	4DCF	19919
x"00",	-- Hex Addr	4DD0	19920
x"00",	-- Hex Addr	4DD1	19921
x"00",	-- Hex Addr	4DD2	19922
x"00",	-- Hex Addr	4DD3	19923
x"00",	-- Hex Addr	4DD4	19924
x"00",	-- Hex Addr	4DD5	19925
x"00",	-- Hex Addr	4DD6	19926
x"00",	-- Hex Addr	4DD7	19927
x"00",	-- Hex Addr	4DD8	19928
x"00",	-- Hex Addr	4DD9	19929
x"00",	-- Hex Addr	4DDA	19930
x"00",	-- Hex Addr	4DDB	19931
x"00",	-- Hex Addr	4DDC	19932
x"00",	-- Hex Addr	4DDD	19933
x"00",	-- Hex Addr	4DDE	19934
x"00",	-- Hex Addr	4DDF	19935
x"00",	-- Hex Addr	4DE0	19936
x"00",	-- Hex Addr	4DE1	19937
x"00",	-- Hex Addr	4DE2	19938
x"00",	-- Hex Addr	4DE3	19939
x"00",	-- Hex Addr	4DE4	19940
x"00",	-- Hex Addr	4DE5	19941
x"00",	-- Hex Addr	4DE6	19942
x"00",	-- Hex Addr	4DE7	19943
x"00",	-- Hex Addr	4DE8	19944
x"00",	-- Hex Addr	4DE9	19945
x"00",	-- Hex Addr	4DEA	19946
x"00",	-- Hex Addr	4DEB	19947
x"00",	-- Hex Addr	4DEC	19948
x"00",	-- Hex Addr	4DED	19949
x"00",	-- Hex Addr	4DEE	19950
x"00",	-- Hex Addr	4DEF	19951
x"00",	-- Hex Addr	4DF0	19952
x"00",	-- Hex Addr	4DF1	19953
x"00",	-- Hex Addr	4DF2	19954
x"00",	-- Hex Addr	4DF3	19955
x"00",	-- Hex Addr	4DF4	19956
x"00",	-- Hex Addr	4DF5	19957
x"00",	-- Hex Addr	4DF6	19958
x"00",	-- Hex Addr	4DF7	19959
x"00",	-- Hex Addr	4DF8	19960
x"00",	-- Hex Addr	4DF9	19961
x"00",	-- Hex Addr	4DFA	19962
x"00",	-- Hex Addr	4DFB	19963
x"00",	-- Hex Addr	4DFC	19964
x"00",	-- Hex Addr	4DFD	19965
x"00",	-- Hex Addr	4DFE	19966
x"00",	-- Hex Addr	4DFF	19967
x"00",	-- Hex Addr	4E00	19968
x"00",	-- Hex Addr	4E01	19969
x"00",	-- Hex Addr	4E02	19970
x"00",	-- Hex Addr	4E03	19971
x"00",	-- Hex Addr	4E04	19972
x"00",	-- Hex Addr	4E05	19973
x"00",	-- Hex Addr	4E06	19974
x"00",	-- Hex Addr	4E07	19975
x"00",	-- Hex Addr	4E08	19976
x"00",	-- Hex Addr	4E09	19977
x"00",	-- Hex Addr	4E0A	19978
x"00",	-- Hex Addr	4E0B	19979
x"00",	-- Hex Addr	4E0C	19980
x"00",	-- Hex Addr	4E0D	19981
x"00",	-- Hex Addr	4E0E	19982
x"00",	-- Hex Addr	4E0F	19983
x"00",	-- Hex Addr	4E10	19984
x"00",	-- Hex Addr	4E11	19985
x"00",	-- Hex Addr	4E12	19986
x"00",	-- Hex Addr	4E13	19987
x"00",	-- Hex Addr	4E14	19988
x"00",	-- Hex Addr	4E15	19989
x"00",	-- Hex Addr	4E16	19990
x"00",	-- Hex Addr	4E17	19991
x"00",	-- Hex Addr	4E18	19992
x"00",	-- Hex Addr	4E19	19993
x"00",	-- Hex Addr	4E1A	19994
x"00",	-- Hex Addr	4E1B	19995
x"00",	-- Hex Addr	4E1C	19996
x"00",	-- Hex Addr	4E1D	19997
x"00",	-- Hex Addr	4E1E	19998
x"00",	-- Hex Addr	4E1F	19999
x"00",	-- Hex Addr	4E20	20000
x"00",	-- Hex Addr	4E21	20001
x"00",	-- Hex Addr	4E22	20002
x"00",	-- Hex Addr	4E23	20003
x"00",	-- Hex Addr	4E24	20004
x"00",	-- Hex Addr	4E25	20005
x"00",	-- Hex Addr	4E26	20006
x"00",	-- Hex Addr	4E27	20007
x"00",	-- Hex Addr	4E28	20008
x"00",	-- Hex Addr	4E29	20009
x"00",	-- Hex Addr	4E2A	20010
x"00",	-- Hex Addr	4E2B	20011
x"00",	-- Hex Addr	4E2C	20012
x"00",	-- Hex Addr	4E2D	20013
x"00",	-- Hex Addr	4E2E	20014
x"00",	-- Hex Addr	4E2F	20015
x"00",	-- Hex Addr	4E30	20016
x"00",	-- Hex Addr	4E31	20017
x"00",	-- Hex Addr	4E32	20018
x"00",	-- Hex Addr	4E33	20019
x"00",	-- Hex Addr	4E34	20020
x"00",	-- Hex Addr	4E35	20021
x"00",	-- Hex Addr	4E36	20022
x"00",	-- Hex Addr	4E37	20023
x"00",	-- Hex Addr	4E38	20024
x"00",	-- Hex Addr	4E39	20025
x"00",	-- Hex Addr	4E3A	20026
x"00",	-- Hex Addr	4E3B	20027
x"00",	-- Hex Addr	4E3C	20028
x"00",	-- Hex Addr	4E3D	20029
x"00",	-- Hex Addr	4E3E	20030
x"00",	-- Hex Addr	4E3F	20031
x"00",	-- Hex Addr	4E40	20032
x"00",	-- Hex Addr	4E41	20033
x"00",	-- Hex Addr	4E42	20034
x"00",	-- Hex Addr	4E43	20035
x"00",	-- Hex Addr	4E44	20036
x"00",	-- Hex Addr	4E45	20037
x"00",	-- Hex Addr	4E46	20038
x"00",	-- Hex Addr	4E47	20039
x"00",	-- Hex Addr	4E48	20040
x"00",	-- Hex Addr	4E49	20041
x"00",	-- Hex Addr	4E4A	20042
x"00",	-- Hex Addr	4E4B	20043
x"00",	-- Hex Addr	4E4C	20044
x"00",	-- Hex Addr	4E4D	20045
x"00",	-- Hex Addr	4E4E	20046
x"00",	-- Hex Addr	4E4F	20047
x"00",	-- Hex Addr	4E50	20048
x"00",	-- Hex Addr	4E51	20049
x"00",	-- Hex Addr	4E52	20050
x"00",	-- Hex Addr	4E53	20051
x"00",	-- Hex Addr	4E54	20052
x"00",	-- Hex Addr	4E55	20053
x"00",	-- Hex Addr	4E56	20054
x"00",	-- Hex Addr	4E57	20055
x"00",	-- Hex Addr	4E58	20056
x"00",	-- Hex Addr	4E59	20057
x"00",	-- Hex Addr	4E5A	20058
x"00",	-- Hex Addr	4E5B	20059
x"00",	-- Hex Addr	4E5C	20060
x"00",	-- Hex Addr	4E5D	20061
x"00",	-- Hex Addr	4E5E	20062
x"00",	-- Hex Addr	4E5F	20063
x"00",	-- Hex Addr	4E60	20064
x"00",	-- Hex Addr	4E61	20065
x"00",	-- Hex Addr	4E62	20066
x"00",	-- Hex Addr	4E63	20067
x"00",	-- Hex Addr	4E64	20068
x"00",	-- Hex Addr	4E65	20069
x"00",	-- Hex Addr	4E66	20070
x"00",	-- Hex Addr	4E67	20071
x"00",	-- Hex Addr	4E68	20072
x"00",	-- Hex Addr	4E69	20073
x"00",	-- Hex Addr	4E6A	20074
x"00",	-- Hex Addr	4E6B	20075
x"00",	-- Hex Addr	4E6C	20076
x"00",	-- Hex Addr	4E6D	20077
x"00",	-- Hex Addr	4E6E	20078
x"00",	-- Hex Addr	4E6F	20079
x"00",	-- Hex Addr	4E70	20080
x"00",	-- Hex Addr	4E71	20081
x"00",	-- Hex Addr	4E72	20082
x"00",	-- Hex Addr	4E73	20083
x"00",	-- Hex Addr	4E74	20084
x"00",	-- Hex Addr	4E75	20085
x"00",	-- Hex Addr	4E76	20086
x"00",	-- Hex Addr	4E77	20087
x"00",	-- Hex Addr	4E78	20088
x"00",	-- Hex Addr	4E79	20089
x"00",	-- Hex Addr	4E7A	20090
x"00",	-- Hex Addr	4E7B	20091
x"00",	-- Hex Addr	4E7C	20092
x"00",	-- Hex Addr	4E7D	20093
x"00",	-- Hex Addr	4E7E	20094
x"00",	-- Hex Addr	4E7F	20095
x"00",	-- Hex Addr	4E80	20096
x"00",	-- Hex Addr	4E81	20097
x"00",	-- Hex Addr	4E82	20098
x"00",	-- Hex Addr	4E83	20099
x"00",	-- Hex Addr	4E84	20100
x"00",	-- Hex Addr	4E85	20101
x"00",	-- Hex Addr	4E86	20102
x"00",	-- Hex Addr	4E87	20103
x"00",	-- Hex Addr	4E88	20104
x"00",	-- Hex Addr	4E89	20105
x"00",	-- Hex Addr	4E8A	20106
x"00",	-- Hex Addr	4E8B	20107
x"00",	-- Hex Addr	4E8C	20108
x"00",	-- Hex Addr	4E8D	20109
x"00",	-- Hex Addr	4E8E	20110
x"00",	-- Hex Addr	4E8F	20111
x"00",	-- Hex Addr	4E90	20112
x"00",	-- Hex Addr	4E91	20113
x"00",	-- Hex Addr	4E92	20114
x"00",	-- Hex Addr	4E93	20115
x"00",	-- Hex Addr	4E94	20116
x"00",	-- Hex Addr	4E95	20117
x"00",	-- Hex Addr	4E96	20118
x"00",	-- Hex Addr	4E97	20119
x"00",	-- Hex Addr	4E98	20120
x"00",	-- Hex Addr	4E99	20121
x"00",	-- Hex Addr	4E9A	20122
x"00",	-- Hex Addr	4E9B	20123
x"00",	-- Hex Addr	4E9C	20124
x"00",	-- Hex Addr	4E9D	20125
x"00",	-- Hex Addr	4E9E	20126
x"00",	-- Hex Addr	4E9F	20127
x"00",	-- Hex Addr	4EA0	20128
x"00",	-- Hex Addr	4EA1	20129
x"00",	-- Hex Addr	4EA2	20130
x"00",	-- Hex Addr	4EA3	20131
x"00",	-- Hex Addr	4EA4	20132
x"00",	-- Hex Addr	4EA5	20133
x"00",	-- Hex Addr	4EA6	20134
x"00",	-- Hex Addr	4EA7	20135
x"00",	-- Hex Addr	4EA8	20136
x"00",	-- Hex Addr	4EA9	20137
x"00",	-- Hex Addr	4EAA	20138
x"00",	-- Hex Addr	4EAB	20139
x"00",	-- Hex Addr	4EAC	20140
x"00",	-- Hex Addr	4EAD	20141
x"00",	-- Hex Addr	4EAE	20142
x"00",	-- Hex Addr	4EAF	20143
x"00",	-- Hex Addr	4EB0	20144
x"00",	-- Hex Addr	4EB1	20145
x"00",	-- Hex Addr	4EB2	20146
x"00",	-- Hex Addr	4EB3	20147
x"00",	-- Hex Addr	4EB4	20148
x"00",	-- Hex Addr	4EB5	20149
x"00",	-- Hex Addr	4EB6	20150
x"00",	-- Hex Addr	4EB7	20151
x"00",	-- Hex Addr	4EB8	20152
x"00",	-- Hex Addr	4EB9	20153
x"00",	-- Hex Addr	4EBA	20154
x"00",	-- Hex Addr	4EBB	20155
x"00",	-- Hex Addr	4EBC	20156
x"00",	-- Hex Addr	4EBD	20157
x"00",	-- Hex Addr	4EBE	20158
x"00",	-- Hex Addr	4EBF	20159
x"00",	-- Hex Addr	4EC0	20160
x"00",	-- Hex Addr	4EC1	20161
x"00",	-- Hex Addr	4EC2	20162
x"00",	-- Hex Addr	4EC3	20163
x"00",	-- Hex Addr	4EC4	20164
x"00",	-- Hex Addr	4EC5	20165
x"00",	-- Hex Addr	4EC6	20166
x"00",	-- Hex Addr	4EC7	20167
x"00",	-- Hex Addr	4EC8	20168
x"00",	-- Hex Addr	4EC9	20169
x"00",	-- Hex Addr	4ECA	20170
x"00",	-- Hex Addr	4ECB	20171
x"00",	-- Hex Addr	4ECC	20172
x"00",	-- Hex Addr	4ECD	20173
x"00",	-- Hex Addr	4ECE	20174
x"00",	-- Hex Addr	4ECF	20175
x"00",	-- Hex Addr	4ED0	20176
x"00",	-- Hex Addr	4ED1	20177
x"00",	-- Hex Addr	4ED2	20178
x"00",	-- Hex Addr	4ED3	20179
x"00",	-- Hex Addr	4ED4	20180
x"00",	-- Hex Addr	4ED5	20181
x"00",	-- Hex Addr	4ED6	20182
x"00",	-- Hex Addr	4ED7	20183
x"00",	-- Hex Addr	4ED8	20184
x"00",	-- Hex Addr	4ED9	20185
x"00",	-- Hex Addr	4EDA	20186
x"00",	-- Hex Addr	4EDB	20187
x"00",	-- Hex Addr	4EDC	20188
x"00",	-- Hex Addr	4EDD	20189
x"00",	-- Hex Addr	4EDE	20190
x"00",	-- Hex Addr	4EDF	20191
x"00",	-- Hex Addr	4EE0	20192
x"00",	-- Hex Addr	4EE1	20193
x"00",	-- Hex Addr	4EE2	20194
x"00",	-- Hex Addr	4EE3	20195
x"00",	-- Hex Addr	4EE4	20196
x"00",	-- Hex Addr	4EE5	20197
x"00",	-- Hex Addr	4EE6	20198
x"00",	-- Hex Addr	4EE7	20199
x"00",	-- Hex Addr	4EE8	20200
x"00",	-- Hex Addr	4EE9	20201
x"00",	-- Hex Addr	4EEA	20202
x"00",	-- Hex Addr	4EEB	20203
x"00",	-- Hex Addr	4EEC	20204
x"00",	-- Hex Addr	4EED	20205
x"00",	-- Hex Addr	4EEE	20206
x"00",	-- Hex Addr	4EEF	20207
x"00",	-- Hex Addr	4EF0	20208
x"00",	-- Hex Addr	4EF1	20209
x"00",	-- Hex Addr	4EF2	20210
x"00",	-- Hex Addr	4EF3	20211
x"00",	-- Hex Addr	4EF4	20212
x"00",	-- Hex Addr	4EF5	20213
x"00",	-- Hex Addr	4EF6	20214
x"00",	-- Hex Addr	4EF7	20215
x"00",	-- Hex Addr	4EF8	20216
x"00",	-- Hex Addr	4EF9	20217
x"00",	-- Hex Addr	4EFA	20218
x"00",	-- Hex Addr	4EFB	20219
x"00",	-- Hex Addr	4EFC	20220
x"00",	-- Hex Addr	4EFD	20221
x"00",	-- Hex Addr	4EFE	20222
x"00",	-- Hex Addr	4EFF	20223
x"00",	-- Hex Addr	4F00	20224
x"00",	-- Hex Addr	4F01	20225
x"00",	-- Hex Addr	4F02	20226
x"00",	-- Hex Addr	4F03	20227
x"00",	-- Hex Addr	4F04	20228
x"00",	-- Hex Addr	4F05	20229
x"00",	-- Hex Addr	4F06	20230
x"00",	-- Hex Addr	4F07	20231
x"00",	-- Hex Addr	4F08	20232
x"00",	-- Hex Addr	4F09	20233
x"00",	-- Hex Addr	4F0A	20234
x"00",	-- Hex Addr	4F0B	20235
x"00",	-- Hex Addr	4F0C	20236
x"00",	-- Hex Addr	4F0D	20237
x"00",	-- Hex Addr	4F0E	20238
x"00",	-- Hex Addr	4F0F	20239
x"00",	-- Hex Addr	4F10	20240
x"00",	-- Hex Addr	4F11	20241
x"00",	-- Hex Addr	4F12	20242
x"00",	-- Hex Addr	4F13	20243
x"00",	-- Hex Addr	4F14	20244
x"00",	-- Hex Addr	4F15	20245
x"00",	-- Hex Addr	4F16	20246
x"00",	-- Hex Addr	4F17	20247
x"00",	-- Hex Addr	4F18	20248
x"00",	-- Hex Addr	4F19	20249
x"00",	-- Hex Addr	4F1A	20250
x"00",	-- Hex Addr	4F1B	20251
x"00",	-- Hex Addr	4F1C	20252
x"00",	-- Hex Addr	4F1D	20253
x"00",	-- Hex Addr	4F1E	20254
x"00",	-- Hex Addr	4F1F	20255
x"00",	-- Hex Addr	4F20	20256
x"00",	-- Hex Addr	4F21	20257
x"00",	-- Hex Addr	4F22	20258
x"00",	-- Hex Addr	4F23	20259
x"00",	-- Hex Addr	4F24	20260
x"00",	-- Hex Addr	4F25	20261
x"00",	-- Hex Addr	4F26	20262
x"00",	-- Hex Addr	4F27	20263
x"00",	-- Hex Addr	4F28	20264
x"00",	-- Hex Addr	4F29	20265
x"00",	-- Hex Addr	4F2A	20266
x"00",	-- Hex Addr	4F2B	20267
x"00",	-- Hex Addr	4F2C	20268
x"00",	-- Hex Addr	4F2D	20269
x"00",	-- Hex Addr	4F2E	20270
x"00",	-- Hex Addr	4F2F	20271
x"00",	-- Hex Addr	4F30	20272
x"00",	-- Hex Addr	4F31	20273
x"00",	-- Hex Addr	4F32	20274
x"00",	-- Hex Addr	4F33	20275
x"00",	-- Hex Addr	4F34	20276
x"00",	-- Hex Addr	4F35	20277
x"00",	-- Hex Addr	4F36	20278
x"00",	-- Hex Addr	4F37	20279
x"00",	-- Hex Addr	4F38	20280
x"00",	-- Hex Addr	4F39	20281
x"00",	-- Hex Addr	4F3A	20282
x"00",	-- Hex Addr	4F3B	20283
x"00",	-- Hex Addr	4F3C	20284
x"00",	-- Hex Addr	4F3D	20285
x"00",	-- Hex Addr	4F3E	20286
x"00",	-- Hex Addr	4F3F	20287
x"00",	-- Hex Addr	4F40	20288
x"00",	-- Hex Addr	4F41	20289
x"00",	-- Hex Addr	4F42	20290
x"00",	-- Hex Addr	4F43	20291
x"00",	-- Hex Addr	4F44	20292
x"00",	-- Hex Addr	4F45	20293
x"00",	-- Hex Addr	4F46	20294
x"00",	-- Hex Addr	4F47	20295
x"00",	-- Hex Addr	4F48	20296
x"00",	-- Hex Addr	4F49	20297
x"00",	-- Hex Addr	4F4A	20298
x"00",	-- Hex Addr	4F4B	20299
x"00",	-- Hex Addr	4F4C	20300
x"00",	-- Hex Addr	4F4D	20301
x"00",	-- Hex Addr	4F4E	20302
x"00",	-- Hex Addr	4F4F	20303
x"00",	-- Hex Addr	4F50	20304
x"00",	-- Hex Addr	4F51	20305
x"00",	-- Hex Addr	4F52	20306
x"00",	-- Hex Addr	4F53	20307
x"00",	-- Hex Addr	4F54	20308
x"00",	-- Hex Addr	4F55	20309
x"00",	-- Hex Addr	4F56	20310
x"00",	-- Hex Addr	4F57	20311
x"00",	-- Hex Addr	4F58	20312
x"00",	-- Hex Addr	4F59	20313
x"00",	-- Hex Addr	4F5A	20314
x"00",	-- Hex Addr	4F5B	20315
x"00",	-- Hex Addr	4F5C	20316
x"00",	-- Hex Addr	4F5D	20317
x"00",	-- Hex Addr	4F5E	20318
x"00",	-- Hex Addr	4F5F	20319
x"00",	-- Hex Addr	4F60	20320
x"00",	-- Hex Addr	4F61	20321
x"00",	-- Hex Addr	4F62	20322
x"00",	-- Hex Addr	4F63	20323
x"00",	-- Hex Addr	4F64	20324
x"00",	-- Hex Addr	4F65	20325
x"00",	-- Hex Addr	4F66	20326
x"00",	-- Hex Addr	4F67	20327
x"00",	-- Hex Addr	4F68	20328
x"00",	-- Hex Addr	4F69	20329
x"00",	-- Hex Addr	4F6A	20330
x"00",	-- Hex Addr	4F6B	20331
x"00",	-- Hex Addr	4F6C	20332
x"00",	-- Hex Addr	4F6D	20333
x"00",	-- Hex Addr	4F6E	20334
x"00",	-- Hex Addr	4F6F	20335
x"00",	-- Hex Addr	4F70	20336
x"00",	-- Hex Addr	4F71	20337
x"00",	-- Hex Addr	4F72	20338
x"00",	-- Hex Addr	4F73	20339
x"00",	-- Hex Addr	4F74	20340
x"00",	-- Hex Addr	4F75	20341
x"00",	-- Hex Addr	4F76	20342
x"00",	-- Hex Addr	4F77	20343
x"00",	-- Hex Addr	4F78	20344
x"00",	-- Hex Addr	4F79	20345
x"00",	-- Hex Addr	4F7A	20346
x"00",	-- Hex Addr	4F7B	20347
x"00",	-- Hex Addr	4F7C	20348
x"00",	-- Hex Addr	4F7D	20349
x"00",	-- Hex Addr	4F7E	20350
x"00",	-- Hex Addr	4F7F	20351
x"00",	-- Hex Addr	4F80	20352
x"00",	-- Hex Addr	4F81	20353
x"00",	-- Hex Addr	4F82	20354
x"00",	-- Hex Addr	4F83	20355
x"00",	-- Hex Addr	4F84	20356
x"00",	-- Hex Addr	4F85	20357
x"00",	-- Hex Addr	4F86	20358
x"00",	-- Hex Addr	4F87	20359
x"00",	-- Hex Addr	4F88	20360
x"00",	-- Hex Addr	4F89	20361
x"00",	-- Hex Addr	4F8A	20362
x"00",	-- Hex Addr	4F8B	20363
x"00",	-- Hex Addr	4F8C	20364
x"00",	-- Hex Addr	4F8D	20365
x"00",	-- Hex Addr	4F8E	20366
x"00",	-- Hex Addr	4F8F	20367
x"00",	-- Hex Addr	4F90	20368
x"00",	-- Hex Addr	4F91	20369
x"00",	-- Hex Addr	4F92	20370
x"00",	-- Hex Addr	4F93	20371
x"00",	-- Hex Addr	4F94	20372
x"00",	-- Hex Addr	4F95	20373
x"00",	-- Hex Addr	4F96	20374
x"00",	-- Hex Addr	4F97	20375
x"00",	-- Hex Addr	4F98	20376
x"00",	-- Hex Addr	4F99	20377
x"00",	-- Hex Addr	4F9A	20378
x"00",	-- Hex Addr	4F9B	20379
x"00",	-- Hex Addr	4F9C	20380
x"00",	-- Hex Addr	4F9D	20381
x"00",	-- Hex Addr	4F9E	20382
x"00",	-- Hex Addr	4F9F	20383
x"00",	-- Hex Addr	4FA0	20384
x"00",	-- Hex Addr	4FA1	20385
x"00",	-- Hex Addr	4FA2	20386
x"00",	-- Hex Addr	4FA3	20387
x"00",	-- Hex Addr	4FA4	20388
x"00",	-- Hex Addr	4FA5	20389
x"00",	-- Hex Addr	4FA6	20390
x"00",	-- Hex Addr	4FA7	20391
x"00",	-- Hex Addr	4FA8	20392
x"00",	-- Hex Addr	4FA9	20393
x"00",	-- Hex Addr	4FAA	20394
x"00",	-- Hex Addr	4FAB	20395
x"00",	-- Hex Addr	4FAC	20396
x"00",	-- Hex Addr	4FAD	20397
x"00",	-- Hex Addr	4FAE	20398
x"00",	-- Hex Addr	4FAF	20399
x"00",	-- Hex Addr	4FB0	20400
x"00",	-- Hex Addr	4FB1	20401
x"00",	-- Hex Addr	4FB2	20402
x"00",	-- Hex Addr	4FB3	20403
x"00",	-- Hex Addr	4FB4	20404
x"00",	-- Hex Addr	4FB5	20405
x"00",	-- Hex Addr	4FB6	20406
x"00",	-- Hex Addr	4FB7	20407
x"00",	-- Hex Addr	4FB8	20408
x"00",	-- Hex Addr	4FB9	20409
x"00",	-- Hex Addr	4FBA	20410
x"00",	-- Hex Addr	4FBB	20411
x"00",	-- Hex Addr	4FBC	20412
x"00",	-- Hex Addr	4FBD	20413
x"00",	-- Hex Addr	4FBE	20414
x"00",	-- Hex Addr	4FBF	20415
x"00",	-- Hex Addr	4FC0	20416
x"00",	-- Hex Addr	4FC1	20417
x"00",	-- Hex Addr	4FC2	20418
x"00",	-- Hex Addr	4FC3	20419
x"00",	-- Hex Addr	4FC4	20420
x"00",	-- Hex Addr	4FC5	20421
x"00",	-- Hex Addr	4FC6	20422
x"00",	-- Hex Addr	4FC7	20423
x"00",	-- Hex Addr	4FC8	20424
x"00",	-- Hex Addr	4FC9	20425
x"00",	-- Hex Addr	4FCA	20426
x"00",	-- Hex Addr	4FCB	20427
x"00",	-- Hex Addr	4FCC	20428
x"00",	-- Hex Addr	4FCD	20429
x"00",	-- Hex Addr	4FCE	20430
x"00",	-- Hex Addr	4FCF	20431
x"00",	-- Hex Addr	4FD0	20432
x"00",	-- Hex Addr	4FD1	20433
x"00",	-- Hex Addr	4FD2	20434
x"00",	-- Hex Addr	4FD3	20435
x"00",	-- Hex Addr	4FD4	20436
x"00",	-- Hex Addr	4FD5	20437
x"00",	-- Hex Addr	4FD6	20438
x"00",	-- Hex Addr	4FD7	20439
x"00",	-- Hex Addr	4FD8	20440
x"00",	-- Hex Addr	4FD9	20441
x"00",	-- Hex Addr	4FDA	20442
x"00",	-- Hex Addr	4FDB	20443
x"00",	-- Hex Addr	4FDC	20444
x"00",	-- Hex Addr	4FDD	20445
x"00",	-- Hex Addr	4FDE	20446
x"00",	-- Hex Addr	4FDF	20447
x"00",	-- Hex Addr	4FE0	20448
x"00",	-- Hex Addr	4FE1	20449
x"00",	-- Hex Addr	4FE2	20450
x"00",	-- Hex Addr	4FE3	20451
x"00",	-- Hex Addr	4FE4	20452
x"00",	-- Hex Addr	4FE5	20453
x"00",	-- Hex Addr	4FE6	20454
x"00",	-- Hex Addr	4FE7	20455
x"00",	-- Hex Addr	4FE8	20456
x"00",	-- Hex Addr	4FE9	20457
x"00",	-- Hex Addr	4FEA	20458
x"00",	-- Hex Addr	4FEB	20459
x"00",	-- Hex Addr	4FEC	20460
x"00",	-- Hex Addr	4FED	20461
x"00",	-- Hex Addr	4FEE	20462
x"00",	-- Hex Addr	4FEF	20463
x"00",	-- Hex Addr	4FF0	20464
x"00",	-- Hex Addr	4FF1	20465
x"00",	-- Hex Addr	4FF2	20466
x"00",	-- Hex Addr	4FF3	20467
x"00",	-- Hex Addr	4FF4	20468
x"00",	-- Hex Addr	4FF5	20469
x"00",	-- Hex Addr	4FF6	20470
x"00",	-- Hex Addr	4FF7	20471
x"00",	-- Hex Addr	4FF8	20472
x"00",	-- Hex Addr	4FF9	20473
x"00",	-- Hex Addr	4FFA	20474
x"00",	-- Hex Addr	4FFB	20475
x"00",	-- Hex Addr	4FFC	20476
x"00",	-- Hex Addr	4FFD	20477
x"00",	-- Hex Addr	4FFE	20478
x"00",	-- Hex Addr	4FFF	20479
x"00",	-- Hex Addr	5000	20480
x"00",	-- Hex Addr	5001	20481
x"00",	-- Hex Addr	5002	20482
x"00",	-- Hex Addr	5003	20483
x"00",	-- Hex Addr	5004	20484
x"00",	-- Hex Addr	5005	20485
x"00",	-- Hex Addr	5006	20486
x"00",	-- Hex Addr	5007	20487
x"00",	-- Hex Addr	5008	20488
x"00",	-- Hex Addr	5009	20489
x"00",	-- Hex Addr	500A	20490
x"00",	-- Hex Addr	500B	20491
x"00",	-- Hex Addr	500C	20492
x"00",	-- Hex Addr	500D	20493
x"00",	-- Hex Addr	500E	20494
x"00",	-- Hex Addr	500F	20495
x"00",	-- Hex Addr	5010	20496
x"00",	-- Hex Addr	5011	20497
x"00",	-- Hex Addr	5012	20498
x"00",	-- Hex Addr	5013	20499
x"00",	-- Hex Addr	5014	20500
x"00",	-- Hex Addr	5015	20501
x"00",	-- Hex Addr	5016	20502
x"00",	-- Hex Addr	5017	20503
x"00",	-- Hex Addr	5018	20504
x"00",	-- Hex Addr	5019	20505
x"00",	-- Hex Addr	501A	20506
x"00",	-- Hex Addr	501B	20507
x"00",	-- Hex Addr	501C	20508
x"00",	-- Hex Addr	501D	20509
x"00",	-- Hex Addr	501E	20510
x"00",	-- Hex Addr	501F	20511
x"00",	-- Hex Addr	5020	20512
x"00",	-- Hex Addr	5021	20513
x"00",	-- Hex Addr	5022	20514
x"00",	-- Hex Addr	5023	20515
x"00",	-- Hex Addr	5024	20516
x"00",	-- Hex Addr	5025	20517
x"00",	-- Hex Addr	5026	20518
x"00",	-- Hex Addr	5027	20519
x"00",	-- Hex Addr	5028	20520
x"00",	-- Hex Addr	5029	20521
x"00",	-- Hex Addr	502A	20522
x"00",	-- Hex Addr	502B	20523
x"00",	-- Hex Addr	502C	20524
x"00",	-- Hex Addr	502D	20525
x"00",	-- Hex Addr	502E	20526
x"00",	-- Hex Addr	502F	20527
x"00",	-- Hex Addr	5030	20528
x"00",	-- Hex Addr	5031	20529
x"00",	-- Hex Addr	5032	20530
x"00",	-- Hex Addr	5033	20531
x"00",	-- Hex Addr	5034	20532
x"00",	-- Hex Addr	5035	20533
x"00",	-- Hex Addr	5036	20534
x"00",	-- Hex Addr	5037	20535
x"00",	-- Hex Addr	5038	20536
x"00",	-- Hex Addr	5039	20537
x"00",	-- Hex Addr	503A	20538
x"00",	-- Hex Addr	503B	20539
x"00",	-- Hex Addr	503C	20540
x"00",	-- Hex Addr	503D	20541
x"00",	-- Hex Addr	503E	20542
x"00",	-- Hex Addr	503F	20543
x"00",	-- Hex Addr	5040	20544
x"00",	-- Hex Addr	5041	20545
x"00",	-- Hex Addr	5042	20546
x"00",	-- Hex Addr	5043	20547
x"00",	-- Hex Addr	5044	20548
x"00",	-- Hex Addr	5045	20549
x"00",	-- Hex Addr	5046	20550
x"00",	-- Hex Addr	5047	20551
x"00",	-- Hex Addr	5048	20552
x"00",	-- Hex Addr	5049	20553
x"00",	-- Hex Addr	504A	20554
x"00",	-- Hex Addr	504B	20555
x"00",	-- Hex Addr	504C	20556
x"00",	-- Hex Addr	504D	20557
x"00",	-- Hex Addr	504E	20558
x"00",	-- Hex Addr	504F	20559
x"00",	-- Hex Addr	5050	20560
x"00",	-- Hex Addr	5051	20561
x"00",	-- Hex Addr	5052	20562
x"00",	-- Hex Addr	5053	20563
x"00",	-- Hex Addr	5054	20564
x"00",	-- Hex Addr	5055	20565
x"00",	-- Hex Addr	5056	20566
x"00",	-- Hex Addr	5057	20567
x"00",	-- Hex Addr	5058	20568
x"00",	-- Hex Addr	5059	20569
x"00",	-- Hex Addr	505A	20570
x"00",	-- Hex Addr	505B	20571
x"00",	-- Hex Addr	505C	20572
x"00",	-- Hex Addr	505D	20573
x"00",	-- Hex Addr	505E	20574
x"00",	-- Hex Addr	505F	20575
x"00",	-- Hex Addr	5060	20576
x"00",	-- Hex Addr	5061	20577
x"00",	-- Hex Addr	5062	20578
x"00",	-- Hex Addr	5063	20579
x"00",	-- Hex Addr	5064	20580
x"00",	-- Hex Addr	5065	20581
x"00",	-- Hex Addr	5066	20582
x"00",	-- Hex Addr	5067	20583
x"00",	-- Hex Addr	5068	20584
x"00",	-- Hex Addr	5069	20585
x"00",	-- Hex Addr	506A	20586
x"00",	-- Hex Addr	506B	20587
x"00",	-- Hex Addr	506C	20588
x"00",	-- Hex Addr	506D	20589
x"00",	-- Hex Addr	506E	20590
x"00",	-- Hex Addr	506F	20591
x"00",	-- Hex Addr	5070	20592
x"00",	-- Hex Addr	5071	20593
x"00",	-- Hex Addr	5072	20594
x"00",	-- Hex Addr	5073	20595
x"00",	-- Hex Addr	5074	20596
x"00",	-- Hex Addr	5075	20597
x"00",	-- Hex Addr	5076	20598
x"00",	-- Hex Addr	5077	20599
x"00",	-- Hex Addr	5078	20600
x"00",	-- Hex Addr	5079	20601
x"00",	-- Hex Addr	507A	20602
x"00",	-- Hex Addr	507B	20603
x"00",	-- Hex Addr	507C	20604
x"00",	-- Hex Addr	507D	20605
x"00",	-- Hex Addr	507E	20606
x"00",	-- Hex Addr	507F	20607
x"00",	-- Hex Addr	5080	20608
x"00",	-- Hex Addr	5081	20609
x"00",	-- Hex Addr	5082	20610
x"00",	-- Hex Addr	5083	20611
x"00",	-- Hex Addr	5084	20612
x"00",	-- Hex Addr	5085	20613
x"00",	-- Hex Addr	5086	20614
x"00",	-- Hex Addr	5087	20615
x"00",	-- Hex Addr	5088	20616
x"00",	-- Hex Addr	5089	20617
x"00",	-- Hex Addr	508A	20618
x"00",	-- Hex Addr	508B	20619
x"00",	-- Hex Addr	508C	20620
x"00",	-- Hex Addr	508D	20621
x"00",	-- Hex Addr	508E	20622
x"00",	-- Hex Addr	508F	20623
x"00",	-- Hex Addr	5090	20624
x"00",	-- Hex Addr	5091	20625
x"00",	-- Hex Addr	5092	20626
x"00",	-- Hex Addr	5093	20627
x"00",	-- Hex Addr	5094	20628
x"00",	-- Hex Addr	5095	20629
x"00",	-- Hex Addr	5096	20630
x"00",	-- Hex Addr	5097	20631
x"00",	-- Hex Addr	5098	20632
x"00",	-- Hex Addr	5099	20633
x"00",	-- Hex Addr	509A	20634
x"00",	-- Hex Addr	509B	20635
x"00",	-- Hex Addr	509C	20636
x"00",	-- Hex Addr	509D	20637
x"00",	-- Hex Addr	509E	20638
x"00",	-- Hex Addr	509F	20639
x"00",	-- Hex Addr	50A0	20640
x"00",	-- Hex Addr	50A1	20641
x"00",	-- Hex Addr	50A2	20642
x"00",	-- Hex Addr	50A3	20643
x"00",	-- Hex Addr	50A4	20644
x"00",	-- Hex Addr	50A5	20645
x"00",	-- Hex Addr	50A6	20646
x"00",	-- Hex Addr	50A7	20647
x"00",	-- Hex Addr	50A8	20648
x"00",	-- Hex Addr	50A9	20649
x"00",	-- Hex Addr	50AA	20650
x"00",	-- Hex Addr	50AB	20651
x"00",	-- Hex Addr	50AC	20652
x"00",	-- Hex Addr	50AD	20653
x"00",	-- Hex Addr	50AE	20654
x"00",	-- Hex Addr	50AF	20655
x"00",	-- Hex Addr	50B0	20656
x"00",	-- Hex Addr	50B1	20657
x"00",	-- Hex Addr	50B2	20658
x"00",	-- Hex Addr	50B3	20659
x"00",	-- Hex Addr	50B4	20660
x"00",	-- Hex Addr	50B5	20661
x"00",	-- Hex Addr	50B6	20662
x"00",	-- Hex Addr	50B7	20663
x"00",	-- Hex Addr	50B8	20664
x"00",	-- Hex Addr	50B9	20665
x"00",	-- Hex Addr	50BA	20666
x"00",	-- Hex Addr	50BB	20667
x"00",	-- Hex Addr	50BC	20668
x"00",	-- Hex Addr	50BD	20669
x"00",	-- Hex Addr	50BE	20670
x"00",	-- Hex Addr	50BF	20671
x"00",	-- Hex Addr	50C0	20672
x"00",	-- Hex Addr	50C1	20673
x"00",	-- Hex Addr	50C2	20674
x"00",	-- Hex Addr	50C3	20675
x"00",	-- Hex Addr	50C4	20676
x"00",	-- Hex Addr	50C5	20677
x"00",	-- Hex Addr	50C6	20678
x"00",	-- Hex Addr	50C7	20679
x"00",	-- Hex Addr	50C8	20680
x"00",	-- Hex Addr	50C9	20681
x"00",	-- Hex Addr	50CA	20682
x"00",	-- Hex Addr	50CB	20683
x"00",	-- Hex Addr	50CC	20684
x"00",	-- Hex Addr	50CD	20685
x"00",	-- Hex Addr	50CE	20686
x"00",	-- Hex Addr	50CF	20687
x"00",	-- Hex Addr	50D0	20688
x"00",	-- Hex Addr	50D1	20689
x"00",	-- Hex Addr	50D2	20690
x"00",	-- Hex Addr	50D3	20691
x"00",	-- Hex Addr	50D4	20692
x"00",	-- Hex Addr	50D5	20693
x"00",	-- Hex Addr	50D6	20694
x"00",	-- Hex Addr	50D7	20695
x"00",	-- Hex Addr	50D8	20696
x"00",	-- Hex Addr	50D9	20697
x"00",	-- Hex Addr	50DA	20698
x"00",	-- Hex Addr	50DB	20699
x"00",	-- Hex Addr	50DC	20700
x"00",	-- Hex Addr	50DD	20701
x"00",	-- Hex Addr	50DE	20702
x"00",	-- Hex Addr	50DF	20703
x"00",	-- Hex Addr	50E0	20704
x"00",	-- Hex Addr	50E1	20705
x"00",	-- Hex Addr	50E2	20706
x"00",	-- Hex Addr	50E3	20707
x"00",	-- Hex Addr	50E4	20708
x"00",	-- Hex Addr	50E5	20709
x"00",	-- Hex Addr	50E6	20710
x"00",	-- Hex Addr	50E7	20711
x"00",	-- Hex Addr	50E8	20712
x"00",	-- Hex Addr	50E9	20713
x"00",	-- Hex Addr	50EA	20714
x"00",	-- Hex Addr	50EB	20715
x"00",	-- Hex Addr	50EC	20716
x"00",	-- Hex Addr	50ED	20717
x"00",	-- Hex Addr	50EE	20718
x"00",	-- Hex Addr	50EF	20719
x"00",	-- Hex Addr	50F0	20720
x"00",	-- Hex Addr	50F1	20721
x"00",	-- Hex Addr	50F2	20722
x"00",	-- Hex Addr	50F3	20723
x"00",	-- Hex Addr	50F4	20724
x"00",	-- Hex Addr	50F5	20725
x"00",	-- Hex Addr	50F6	20726
x"00",	-- Hex Addr	50F7	20727
x"00",	-- Hex Addr	50F8	20728
x"00",	-- Hex Addr	50F9	20729
x"00",	-- Hex Addr	50FA	20730
x"00",	-- Hex Addr	50FB	20731
x"00",	-- Hex Addr	50FC	20732
x"00",	-- Hex Addr	50FD	20733
x"00",	-- Hex Addr	50FE	20734
x"00",	-- Hex Addr	50FF	20735
x"00",	-- Hex Addr	5100	20736
x"00",	-- Hex Addr	5101	20737
x"00",	-- Hex Addr	5102	20738
x"00",	-- Hex Addr	5103	20739
x"00",	-- Hex Addr	5104	20740
x"00",	-- Hex Addr	5105	20741
x"00",	-- Hex Addr	5106	20742
x"00",	-- Hex Addr	5107	20743
x"00",	-- Hex Addr	5108	20744
x"00",	-- Hex Addr	5109	20745
x"00",	-- Hex Addr	510A	20746
x"00",	-- Hex Addr	510B	20747
x"00",	-- Hex Addr	510C	20748
x"00",	-- Hex Addr	510D	20749
x"00",	-- Hex Addr	510E	20750
x"00",	-- Hex Addr	510F	20751
x"00",	-- Hex Addr	5110	20752
x"00",	-- Hex Addr	5111	20753
x"00",	-- Hex Addr	5112	20754
x"00",	-- Hex Addr	5113	20755
x"00",	-- Hex Addr	5114	20756
x"00",	-- Hex Addr	5115	20757
x"00",	-- Hex Addr	5116	20758
x"00",	-- Hex Addr	5117	20759
x"00",	-- Hex Addr	5118	20760
x"00",	-- Hex Addr	5119	20761
x"00",	-- Hex Addr	511A	20762
x"00",	-- Hex Addr	511B	20763
x"00",	-- Hex Addr	511C	20764
x"00",	-- Hex Addr	511D	20765
x"00",	-- Hex Addr	511E	20766
x"00",	-- Hex Addr	511F	20767
x"00",	-- Hex Addr	5120	20768
x"00",	-- Hex Addr	5121	20769
x"00",	-- Hex Addr	5122	20770
x"00",	-- Hex Addr	5123	20771
x"00",	-- Hex Addr	5124	20772
x"00",	-- Hex Addr	5125	20773
x"00",	-- Hex Addr	5126	20774
x"00",	-- Hex Addr	5127	20775
x"00",	-- Hex Addr	5128	20776
x"00",	-- Hex Addr	5129	20777
x"00",	-- Hex Addr	512A	20778
x"00",	-- Hex Addr	512B	20779
x"00",	-- Hex Addr	512C	20780
x"00",	-- Hex Addr	512D	20781
x"00",	-- Hex Addr	512E	20782
x"00",	-- Hex Addr	512F	20783
x"00",	-- Hex Addr	5130	20784
x"00",	-- Hex Addr	5131	20785
x"00",	-- Hex Addr	5132	20786
x"00",	-- Hex Addr	5133	20787
x"00",	-- Hex Addr	5134	20788
x"00",	-- Hex Addr	5135	20789
x"00",	-- Hex Addr	5136	20790
x"00",	-- Hex Addr	5137	20791
x"00",	-- Hex Addr	5138	20792
x"00",	-- Hex Addr	5139	20793
x"00",	-- Hex Addr	513A	20794
x"00",	-- Hex Addr	513B	20795
x"00",	-- Hex Addr	513C	20796
x"00",	-- Hex Addr	513D	20797
x"00",	-- Hex Addr	513E	20798
x"00",	-- Hex Addr	513F	20799
x"00",	-- Hex Addr	5140	20800
x"00",	-- Hex Addr	5141	20801
x"00",	-- Hex Addr	5142	20802
x"00",	-- Hex Addr	5143	20803
x"00",	-- Hex Addr	5144	20804
x"00",	-- Hex Addr	5145	20805
x"00",	-- Hex Addr	5146	20806
x"00",	-- Hex Addr	5147	20807
x"00",	-- Hex Addr	5148	20808
x"00",	-- Hex Addr	5149	20809
x"00",	-- Hex Addr	514A	20810
x"00",	-- Hex Addr	514B	20811
x"00",	-- Hex Addr	514C	20812
x"00",	-- Hex Addr	514D	20813
x"00",	-- Hex Addr	514E	20814
x"00",	-- Hex Addr	514F	20815
x"00",	-- Hex Addr	5150	20816
x"00",	-- Hex Addr	5151	20817
x"00",	-- Hex Addr	5152	20818
x"00",	-- Hex Addr	5153	20819
x"00",	-- Hex Addr	5154	20820
x"00",	-- Hex Addr	5155	20821
x"00",	-- Hex Addr	5156	20822
x"00",	-- Hex Addr	5157	20823
x"00",	-- Hex Addr	5158	20824
x"00",	-- Hex Addr	5159	20825
x"00",	-- Hex Addr	515A	20826
x"00",	-- Hex Addr	515B	20827
x"00",	-- Hex Addr	515C	20828
x"00",	-- Hex Addr	515D	20829
x"00",	-- Hex Addr	515E	20830
x"00",	-- Hex Addr	515F	20831
x"00",	-- Hex Addr	5160	20832
x"00",	-- Hex Addr	5161	20833
x"00",	-- Hex Addr	5162	20834
x"00",	-- Hex Addr	5163	20835
x"00",	-- Hex Addr	5164	20836
x"00",	-- Hex Addr	5165	20837
x"00",	-- Hex Addr	5166	20838
x"00",	-- Hex Addr	5167	20839
x"00",	-- Hex Addr	5168	20840
x"00",	-- Hex Addr	5169	20841
x"00",	-- Hex Addr	516A	20842
x"00",	-- Hex Addr	516B	20843
x"00",	-- Hex Addr	516C	20844
x"00",	-- Hex Addr	516D	20845
x"00",	-- Hex Addr	516E	20846
x"00",	-- Hex Addr	516F	20847
x"00",	-- Hex Addr	5170	20848
x"00",	-- Hex Addr	5171	20849
x"00",	-- Hex Addr	5172	20850
x"00",	-- Hex Addr	5173	20851
x"00",	-- Hex Addr	5174	20852
x"00",	-- Hex Addr	5175	20853
x"00",	-- Hex Addr	5176	20854
x"00",	-- Hex Addr	5177	20855
x"00",	-- Hex Addr	5178	20856
x"00",	-- Hex Addr	5179	20857
x"00",	-- Hex Addr	517A	20858
x"00",	-- Hex Addr	517B	20859
x"00",	-- Hex Addr	517C	20860
x"00",	-- Hex Addr	517D	20861
x"00",	-- Hex Addr	517E	20862
x"00",	-- Hex Addr	517F	20863
x"00",	-- Hex Addr	5180	20864
x"00",	-- Hex Addr	5181	20865
x"00",	-- Hex Addr	5182	20866
x"00",	-- Hex Addr	5183	20867
x"00",	-- Hex Addr	5184	20868
x"00",	-- Hex Addr	5185	20869
x"00",	-- Hex Addr	5186	20870
x"00",	-- Hex Addr	5187	20871
x"00",	-- Hex Addr	5188	20872
x"00",	-- Hex Addr	5189	20873
x"00",	-- Hex Addr	518A	20874
x"00",	-- Hex Addr	518B	20875
x"00",	-- Hex Addr	518C	20876
x"00",	-- Hex Addr	518D	20877
x"00",	-- Hex Addr	518E	20878
x"00",	-- Hex Addr	518F	20879
x"00",	-- Hex Addr	5190	20880
x"00",	-- Hex Addr	5191	20881
x"00",	-- Hex Addr	5192	20882
x"00",	-- Hex Addr	5193	20883
x"00",	-- Hex Addr	5194	20884
x"00",	-- Hex Addr	5195	20885
x"00",	-- Hex Addr	5196	20886
x"00",	-- Hex Addr	5197	20887
x"00",	-- Hex Addr	5198	20888
x"00",	-- Hex Addr	5199	20889
x"00",	-- Hex Addr	519A	20890
x"00",	-- Hex Addr	519B	20891
x"00",	-- Hex Addr	519C	20892
x"00",	-- Hex Addr	519D	20893
x"00",	-- Hex Addr	519E	20894
x"00",	-- Hex Addr	519F	20895
x"00",	-- Hex Addr	51A0	20896
x"00",	-- Hex Addr	51A1	20897
x"00",	-- Hex Addr	51A2	20898
x"00",	-- Hex Addr	51A3	20899
x"00",	-- Hex Addr	51A4	20900
x"00",	-- Hex Addr	51A5	20901
x"00",	-- Hex Addr	51A6	20902
x"00",	-- Hex Addr	51A7	20903
x"00",	-- Hex Addr	51A8	20904
x"00",	-- Hex Addr	51A9	20905
x"00",	-- Hex Addr	51AA	20906
x"00",	-- Hex Addr	51AB	20907
x"00",	-- Hex Addr	51AC	20908
x"00",	-- Hex Addr	51AD	20909
x"00",	-- Hex Addr	51AE	20910
x"00",	-- Hex Addr	51AF	20911
x"00",	-- Hex Addr	51B0	20912
x"00",	-- Hex Addr	51B1	20913
x"00",	-- Hex Addr	51B2	20914
x"00",	-- Hex Addr	51B3	20915
x"00",	-- Hex Addr	51B4	20916
x"00",	-- Hex Addr	51B5	20917
x"00",	-- Hex Addr	51B6	20918
x"00",	-- Hex Addr	51B7	20919
x"00",	-- Hex Addr	51B8	20920
x"00",	-- Hex Addr	51B9	20921
x"00",	-- Hex Addr	51BA	20922
x"00",	-- Hex Addr	51BB	20923
x"00",	-- Hex Addr	51BC	20924
x"00",	-- Hex Addr	51BD	20925
x"00",	-- Hex Addr	51BE	20926
x"00",	-- Hex Addr	51BF	20927
x"00",	-- Hex Addr	51C0	20928
x"00",	-- Hex Addr	51C1	20929
x"00",	-- Hex Addr	51C2	20930
x"00",	-- Hex Addr	51C3	20931
x"00",	-- Hex Addr	51C4	20932
x"00",	-- Hex Addr	51C5	20933
x"00",	-- Hex Addr	51C6	20934
x"00",	-- Hex Addr	51C7	20935
x"00",	-- Hex Addr	51C8	20936
x"00",	-- Hex Addr	51C9	20937
x"00",	-- Hex Addr	51CA	20938
x"00",	-- Hex Addr	51CB	20939
x"00",	-- Hex Addr	51CC	20940
x"00",	-- Hex Addr	51CD	20941
x"00",	-- Hex Addr	51CE	20942
x"00",	-- Hex Addr	51CF	20943
x"00",	-- Hex Addr	51D0	20944
x"00",	-- Hex Addr	51D1	20945
x"00",	-- Hex Addr	51D2	20946
x"00",	-- Hex Addr	51D3	20947
x"00",	-- Hex Addr	51D4	20948
x"00",	-- Hex Addr	51D5	20949
x"00",	-- Hex Addr	51D6	20950
x"00",	-- Hex Addr	51D7	20951
x"00",	-- Hex Addr	51D8	20952
x"00",	-- Hex Addr	51D9	20953
x"00",	-- Hex Addr	51DA	20954
x"00",	-- Hex Addr	51DB	20955
x"00",	-- Hex Addr	51DC	20956
x"00",	-- Hex Addr	51DD	20957
x"00",	-- Hex Addr	51DE	20958
x"00",	-- Hex Addr	51DF	20959
x"00",	-- Hex Addr	51E0	20960
x"00",	-- Hex Addr	51E1	20961
x"00",	-- Hex Addr	51E2	20962
x"00",	-- Hex Addr	51E3	20963
x"00",	-- Hex Addr	51E4	20964
x"00",	-- Hex Addr	51E5	20965
x"00",	-- Hex Addr	51E6	20966
x"00",	-- Hex Addr	51E7	20967
x"00",	-- Hex Addr	51E8	20968
x"00",	-- Hex Addr	51E9	20969
x"00",	-- Hex Addr	51EA	20970
x"00",	-- Hex Addr	51EB	20971
x"00",	-- Hex Addr	51EC	20972
x"00",	-- Hex Addr	51ED	20973
x"00",	-- Hex Addr	51EE	20974
x"00",	-- Hex Addr	51EF	20975
x"00",	-- Hex Addr	51F0	20976
x"00",	-- Hex Addr	51F1	20977
x"00",	-- Hex Addr	51F2	20978
x"00",	-- Hex Addr	51F3	20979
x"00",	-- Hex Addr	51F4	20980
x"00",	-- Hex Addr	51F5	20981
x"00",	-- Hex Addr	51F6	20982
x"00",	-- Hex Addr	51F7	20983
x"00",	-- Hex Addr	51F8	20984
x"00",	-- Hex Addr	51F9	20985
x"00",	-- Hex Addr	51FA	20986
x"00",	-- Hex Addr	51FB	20987
x"00",	-- Hex Addr	51FC	20988
x"00",	-- Hex Addr	51FD	20989
x"00",	-- Hex Addr	51FE	20990
x"00",	-- Hex Addr	51FF	20991
x"00",	-- Hex Addr	5200	20992
x"00",	-- Hex Addr	5201	20993
x"00",	-- Hex Addr	5202	20994
x"00",	-- Hex Addr	5203	20995
x"00",	-- Hex Addr	5204	20996
x"00",	-- Hex Addr	5205	20997
x"00",	-- Hex Addr	5206	20998
x"00",	-- Hex Addr	5207	20999
x"00",	-- Hex Addr	5208	21000
x"00",	-- Hex Addr	5209	21001
x"00",	-- Hex Addr	520A	21002
x"00",	-- Hex Addr	520B	21003
x"00",	-- Hex Addr	520C	21004
x"00",	-- Hex Addr	520D	21005
x"00",	-- Hex Addr	520E	21006
x"00",	-- Hex Addr	520F	21007
x"00",	-- Hex Addr	5210	21008
x"00",	-- Hex Addr	5211	21009
x"00",	-- Hex Addr	5212	21010
x"00",	-- Hex Addr	5213	21011
x"00",	-- Hex Addr	5214	21012
x"00",	-- Hex Addr	5215	21013
x"00",	-- Hex Addr	5216	21014
x"00",	-- Hex Addr	5217	21015
x"00",	-- Hex Addr	5218	21016
x"00",	-- Hex Addr	5219	21017
x"00",	-- Hex Addr	521A	21018
x"00",	-- Hex Addr	521B	21019
x"00",	-- Hex Addr	521C	21020
x"00",	-- Hex Addr	521D	21021
x"00",	-- Hex Addr	521E	21022
x"00",	-- Hex Addr	521F	21023
x"00",	-- Hex Addr	5220	21024
x"00",	-- Hex Addr	5221	21025
x"00",	-- Hex Addr	5222	21026
x"00",	-- Hex Addr	5223	21027
x"00",	-- Hex Addr	5224	21028
x"00",	-- Hex Addr	5225	21029
x"00",	-- Hex Addr	5226	21030
x"00",	-- Hex Addr	5227	21031
x"00",	-- Hex Addr	5228	21032
x"00",	-- Hex Addr	5229	21033
x"00",	-- Hex Addr	522A	21034
x"00",	-- Hex Addr	522B	21035
x"00",	-- Hex Addr	522C	21036
x"00",	-- Hex Addr	522D	21037
x"00",	-- Hex Addr	522E	21038
x"00",	-- Hex Addr	522F	21039
x"00",	-- Hex Addr	5230	21040
x"00",	-- Hex Addr	5231	21041
x"00",	-- Hex Addr	5232	21042
x"00",	-- Hex Addr	5233	21043
x"00",	-- Hex Addr	5234	21044
x"00",	-- Hex Addr	5235	21045
x"00",	-- Hex Addr	5236	21046
x"00",	-- Hex Addr	5237	21047
x"00",	-- Hex Addr	5238	21048
x"00",	-- Hex Addr	5239	21049
x"00",	-- Hex Addr	523A	21050
x"00",	-- Hex Addr	523B	21051
x"00",	-- Hex Addr	523C	21052
x"00",	-- Hex Addr	523D	21053
x"00",	-- Hex Addr	523E	21054
x"00",	-- Hex Addr	523F	21055
x"00",	-- Hex Addr	5240	21056
x"00",	-- Hex Addr	5241	21057
x"00",	-- Hex Addr	5242	21058
x"00",	-- Hex Addr	5243	21059
x"00",	-- Hex Addr	5244	21060
x"00",	-- Hex Addr	5245	21061
x"00",	-- Hex Addr	5246	21062
x"00",	-- Hex Addr	5247	21063
x"00",	-- Hex Addr	5248	21064
x"00",	-- Hex Addr	5249	21065
x"00",	-- Hex Addr	524A	21066
x"00",	-- Hex Addr	524B	21067
x"00",	-- Hex Addr	524C	21068
x"00",	-- Hex Addr	524D	21069
x"00",	-- Hex Addr	524E	21070
x"00",	-- Hex Addr	524F	21071
x"00",	-- Hex Addr	5250	21072
x"00",	-- Hex Addr	5251	21073
x"00",	-- Hex Addr	5252	21074
x"00",	-- Hex Addr	5253	21075
x"00",	-- Hex Addr	5254	21076
x"00",	-- Hex Addr	5255	21077
x"00",	-- Hex Addr	5256	21078
x"00",	-- Hex Addr	5257	21079
x"00",	-- Hex Addr	5258	21080
x"00",	-- Hex Addr	5259	21081
x"00",	-- Hex Addr	525A	21082
x"00",	-- Hex Addr	525B	21083
x"00",	-- Hex Addr	525C	21084
x"00",	-- Hex Addr	525D	21085
x"00",	-- Hex Addr	525E	21086
x"00",	-- Hex Addr	525F	21087
x"00",	-- Hex Addr	5260	21088
x"00",	-- Hex Addr	5261	21089
x"00",	-- Hex Addr	5262	21090
x"00",	-- Hex Addr	5263	21091
x"00",	-- Hex Addr	5264	21092
x"00",	-- Hex Addr	5265	21093
x"00",	-- Hex Addr	5266	21094
x"00",	-- Hex Addr	5267	21095
x"00",	-- Hex Addr	5268	21096
x"00",	-- Hex Addr	5269	21097
x"00",	-- Hex Addr	526A	21098
x"00",	-- Hex Addr	526B	21099
x"00",	-- Hex Addr	526C	21100
x"00",	-- Hex Addr	526D	21101
x"00",	-- Hex Addr	526E	21102
x"00",	-- Hex Addr	526F	21103
x"00",	-- Hex Addr	5270	21104
x"00",	-- Hex Addr	5271	21105
x"00",	-- Hex Addr	5272	21106
x"00",	-- Hex Addr	5273	21107
x"00",	-- Hex Addr	5274	21108
x"00",	-- Hex Addr	5275	21109
x"00",	-- Hex Addr	5276	21110
x"00",	-- Hex Addr	5277	21111
x"00",	-- Hex Addr	5278	21112
x"00",	-- Hex Addr	5279	21113
x"00",	-- Hex Addr	527A	21114
x"00",	-- Hex Addr	527B	21115
x"00",	-- Hex Addr	527C	21116
x"00",	-- Hex Addr	527D	21117
x"00",	-- Hex Addr	527E	21118
x"00",	-- Hex Addr	527F	21119
x"00",	-- Hex Addr	5280	21120
x"00",	-- Hex Addr	5281	21121
x"00",	-- Hex Addr	5282	21122
x"00",	-- Hex Addr	5283	21123
x"00",	-- Hex Addr	5284	21124
x"00",	-- Hex Addr	5285	21125
x"00",	-- Hex Addr	5286	21126
x"00",	-- Hex Addr	5287	21127
x"00",	-- Hex Addr	5288	21128
x"00",	-- Hex Addr	5289	21129
x"00",	-- Hex Addr	528A	21130
x"00",	-- Hex Addr	528B	21131
x"00",	-- Hex Addr	528C	21132
x"00",	-- Hex Addr	528D	21133
x"00",	-- Hex Addr	528E	21134
x"00",	-- Hex Addr	528F	21135
x"00",	-- Hex Addr	5290	21136
x"00",	-- Hex Addr	5291	21137
x"00",	-- Hex Addr	5292	21138
x"00",	-- Hex Addr	5293	21139
x"00",	-- Hex Addr	5294	21140
x"00",	-- Hex Addr	5295	21141
x"00",	-- Hex Addr	5296	21142
x"00",	-- Hex Addr	5297	21143
x"00",	-- Hex Addr	5298	21144
x"00",	-- Hex Addr	5299	21145
x"00",	-- Hex Addr	529A	21146
x"00",	-- Hex Addr	529B	21147
x"00",	-- Hex Addr	529C	21148
x"00",	-- Hex Addr	529D	21149
x"00",	-- Hex Addr	529E	21150
x"00",	-- Hex Addr	529F	21151
x"00",	-- Hex Addr	52A0	21152
x"00",	-- Hex Addr	52A1	21153
x"00",	-- Hex Addr	52A2	21154
x"00",	-- Hex Addr	52A3	21155
x"00",	-- Hex Addr	52A4	21156
x"00",	-- Hex Addr	52A5	21157
x"00",	-- Hex Addr	52A6	21158
x"00",	-- Hex Addr	52A7	21159
x"00",	-- Hex Addr	52A8	21160
x"00",	-- Hex Addr	52A9	21161
x"00",	-- Hex Addr	52AA	21162
x"00",	-- Hex Addr	52AB	21163
x"00",	-- Hex Addr	52AC	21164
x"00",	-- Hex Addr	52AD	21165
x"00",	-- Hex Addr	52AE	21166
x"00",	-- Hex Addr	52AF	21167
x"00",	-- Hex Addr	52B0	21168
x"00",	-- Hex Addr	52B1	21169
x"00",	-- Hex Addr	52B2	21170
x"00",	-- Hex Addr	52B3	21171
x"00",	-- Hex Addr	52B4	21172
x"00",	-- Hex Addr	52B5	21173
x"00",	-- Hex Addr	52B6	21174
x"00",	-- Hex Addr	52B7	21175
x"00",	-- Hex Addr	52B8	21176
x"00",	-- Hex Addr	52B9	21177
x"00",	-- Hex Addr	52BA	21178
x"00",	-- Hex Addr	52BB	21179
x"00",	-- Hex Addr	52BC	21180
x"00",	-- Hex Addr	52BD	21181
x"00",	-- Hex Addr	52BE	21182
x"00",	-- Hex Addr	52BF	21183
x"00",	-- Hex Addr	52C0	21184
x"00",	-- Hex Addr	52C1	21185
x"00",	-- Hex Addr	52C2	21186
x"00",	-- Hex Addr	52C3	21187
x"00",	-- Hex Addr	52C4	21188
x"00",	-- Hex Addr	52C5	21189
x"00",	-- Hex Addr	52C6	21190
x"00",	-- Hex Addr	52C7	21191
x"00",	-- Hex Addr	52C8	21192
x"00",	-- Hex Addr	52C9	21193
x"00",	-- Hex Addr	52CA	21194
x"00",	-- Hex Addr	52CB	21195
x"00",	-- Hex Addr	52CC	21196
x"00",	-- Hex Addr	52CD	21197
x"00",	-- Hex Addr	52CE	21198
x"00",	-- Hex Addr	52CF	21199
x"00",	-- Hex Addr	52D0	21200
x"00",	-- Hex Addr	52D1	21201
x"00",	-- Hex Addr	52D2	21202
x"00",	-- Hex Addr	52D3	21203
x"00",	-- Hex Addr	52D4	21204
x"00",	-- Hex Addr	52D5	21205
x"00",	-- Hex Addr	52D6	21206
x"00",	-- Hex Addr	52D7	21207
x"00",	-- Hex Addr	52D8	21208
x"00",	-- Hex Addr	52D9	21209
x"00",	-- Hex Addr	52DA	21210
x"00",	-- Hex Addr	52DB	21211
x"00",	-- Hex Addr	52DC	21212
x"00",	-- Hex Addr	52DD	21213
x"00",	-- Hex Addr	52DE	21214
x"00",	-- Hex Addr	52DF	21215
x"00",	-- Hex Addr	52E0	21216
x"00",	-- Hex Addr	52E1	21217
x"00",	-- Hex Addr	52E2	21218
x"00",	-- Hex Addr	52E3	21219
x"00",	-- Hex Addr	52E4	21220
x"00",	-- Hex Addr	52E5	21221
x"00",	-- Hex Addr	52E6	21222
x"00",	-- Hex Addr	52E7	21223
x"00",	-- Hex Addr	52E8	21224
x"00",	-- Hex Addr	52E9	21225
x"00",	-- Hex Addr	52EA	21226
x"00",	-- Hex Addr	52EB	21227
x"00",	-- Hex Addr	52EC	21228
x"00",	-- Hex Addr	52ED	21229
x"00",	-- Hex Addr	52EE	21230
x"00",	-- Hex Addr	52EF	21231
x"00",	-- Hex Addr	52F0	21232
x"00",	-- Hex Addr	52F1	21233
x"00",	-- Hex Addr	52F2	21234
x"00",	-- Hex Addr	52F3	21235
x"00",	-- Hex Addr	52F4	21236
x"00",	-- Hex Addr	52F5	21237
x"00",	-- Hex Addr	52F6	21238
x"00",	-- Hex Addr	52F7	21239
x"00",	-- Hex Addr	52F8	21240
x"00",	-- Hex Addr	52F9	21241
x"00",	-- Hex Addr	52FA	21242
x"00",	-- Hex Addr	52FB	21243
x"00",	-- Hex Addr	52FC	21244
x"00",	-- Hex Addr	52FD	21245
x"00",	-- Hex Addr	52FE	21246
x"00",	-- Hex Addr	52FF	21247
x"00",	-- Hex Addr	5300	21248
x"00",	-- Hex Addr	5301	21249
x"00",	-- Hex Addr	5302	21250
x"00",	-- Hex Addr	5303	21251
x"00",	-- Hex Addr	5304	21252
x"00",	-- Hex Addr	5305	21253
x"00",	-- Hex Addr	5306	21254
x"00",	-- Hex Addr	5307	21255
x"00",	-- Hex Addr	5308	21256
x"00",	-- Hex Addr	5309	21257
x"00",	-- Hex Addr	530A	21258
x"00",	-- Hex Addr	530B	21259
x"00",	-- Hex Addr	530C	21260
x"00",	-- Hex Addr	530D	21261
x"00",	-- Hex Addr	530E	21262
x"00",	-- Hex Addr	530F	21263
x"00",	-- Hex Addr	5310	21264
x"00",	-- Hex Addr	5311	21265
x"00",	-- Hex Addr	5312	21266
x"00",	-- Hex Addr	5313	21267
x"00",	-- Hex Addr	5314	21268
x"00",	-- Hex Addr	5315	21269
x"00",	-- Hex Addr	5316	21270
x"00",	-- Hex Addr	5317	21271
x"00",	-- Hex Addr	5318	21272
x"00",	-- Hex Addr	5319	21273
x"00",	-- Hex Addr	531A	21274
x"00",	-- Hex Addr	531B	21275
x"00",	-- Hex Addr	531C	21276
x"00",	-- Hex Addr	531D	21277
x"00",	-- Hex Addr	531E	21278
x"00",	-- Hex Addr	531F	21279
x"00",	-- Hex Addr	5320	21280
x"00",	-- Hex Addr	5321	21281
x"00",	-- Hex Addr	5322	21282
x"00",	-- Hex Addr	5323	21283
x"00",	-- Hex Addr	5324	21284
x"00",	-- Hex Addr	5325	21285
x"00",	-- Hex Addr	5326	21286
x"00",	-- Hex Addr	5327	21287
x"00",	-- Hex Addr	5328	21288
x"00",	-- Hex Addr	5329	21289
x"00",	-- Hex Addr	532A	21290
x"00",	-- Hex Addr	532B	21291
x"00",	-- Hex Addr	532C	21292
x"00",	-- Hex Addr	532D	21293
x"00",	-- Hex Addr	532E	21294
x"00",	-- Hex Addr	532F	21295
x"00",	-- Hex Addr	5330	21296
x"00",	-- Hex Addr	5331	21297
x"00",	-- Hex Addr	5332	21298
x"00",	-- Hex Addr	5333	21299
x"00",	-- Hex Addr	5334	21300
x"00",	-- Hex Addr	5335	21301
x"00",	-- Hex Addr	5336	21302
x"00",	-- Hex Addr	5337	21303
x"00",	-- Hex Addr	5338	21304
x"00",	-- Hex Addr	5339	21305
x"00",	-- Hex Addr	533A	21306
x"00",	-- Hex Addr	533B	21307
x"00",	-- Hex Addr	533C	21308
x"00",	-- Hex Addr	533D	21309
x"00",	-- Hex Addr	533E	21310
x"00",	-- Hex Addr	533F	21311
x"00",	-- Hex Addr	5340	21312
x"00",	-- Hex Addr	5341	21313
x"00",	-- Hex Addr	5342	21314
x"00",	-- Hex Addr	5343	21315
x"00",	-- Hex Addr	5344	21316
x"00",	-- Hex Addr	5345	21317
x"00",	-- Hex Addr	5346	21318
x"00",	-- Hex Addr	5347	21319
x"00",	-- Hex Addr	5348	21320
x"00",	-- Hex Addr	5349	21321
x"00",	-- Hex Addr	534A	21322
x"00",	-- Hex Addr	534B	21323
x"00",	-- Hex Addr	534C	21324
x"00",	-- Hex Addr	534D	21325
x"00",	-- Hex Addr	534E	21326
x"00",	-- Hex Addr	534F	21327
x"00",	-- Hex Addr	5350	21328
x"00",	-- Hex Addr	5351	21329
x"00",	-- Hex Addr	5352	21330
x"00",	-- Hex Addr	5353	21331
x"00",	-- Hex Addr	5354	21332
x"00",	-- Hex Addr	5355	21333
x"00",	-- Hex Addr	5356	21334
x"00",	-- Hex Addr	5357	21335
x"00",	-- Hex Addr	5358	21336
x"00",	-- Hex Addr	5359	21337
x"00",	-- Hex Addr	535A	21338
x"00",	-- Hex Addr	535B	21339
x"00",	-- Hex Addr	535C	21340
x"00",	-- Hex Addr	535D	21341
x"00",	-- Hex Addr	535E	21342
x"00",	-- Hex Addr	535F	21343
x"00",	-- Hex Addr	5360	21344
x"00",	-- Hex Addr	5361	21345
x"00",	-- Hex Addr	5362	21346
x"00",	-- Hex Addr	5363	21347
x"00",	-- Hex Addr	5364	21348
x"00",	-- Hex Addr	5365	21349
x"00",	-- Hex Addr	5366	21350
x"00",	-- Hex Addr	5367	21351
x"00",	-- Hex Addr	5368	21352
x"00",	-- Hex Addr	5369	21353
x"00",	-- Hex Addr	536A	21354
x"00",	-- Hex Addr	536B	21355
x"00",	-- Hex Addr	536C	21356
x"00",	-- Hex Addr	536D	21357
x"00",	-- Hex Addr	536E	21358
x"00",	-- Hex Addr	536F	21359
x"00",	-- Hex Addr	5370	21360
x"00",	-- Hex Addr	5371	21361
x"00",	-- Hex Addr	5372	21362
x"00",	-- Hex Addr	5373	21363
x"00",	-- Hex Addr	5374	21364
x"00",	-- Hex Addr	5375	21365
x"00",	-- Hex Addr	5376	21366
x"00",	-- Hex Addr	5377	21367
x"00",	-- Hex Addr	5378	21368
x"00",	-- Hex Addr	5379	21369
x"00",	-- Hex Addr	537A	21370
x"00",	-- Hex Addr	537B	21371
x"00",	-- Hex Addr	537C	21372
x"00",	-- Hex Addr	537D	21373
x"00",	-- Hex Addr	537E	21374
x"00",	-- Hex Addr	537F	21375
x"00",	-- Hex Addr	5380	21376
x"00",	-- Hex Addr	5381	21377
x"00",	-- Hex Addr	5382	21378
x"00",	-- Hex Addr	5383	21379
x"00",	-- Hex Addr	5384	21380
x"00",	-- Hex Addr	5385	21381
x"00",	-- Hex Addr	5386	21382
x"00",	-- Hex Addr	5387	21383
x"00",	-- Hex Addr	5388	21384
x"00",	-- Hex Addr	5389	21385
x"00",	-- Hex Addr	538A	21386
x"00",	-- Hex Addr	538B	21387
x"00",	-- Hex Addr	538C	21388
x"00",	-- Hex Addr	538D	21389
x"00",	-- Hex Addr	538E	21390
x"00",	-- Hex Addr	538F	21391
x"00",	-- Hex Addr	5390	21392
x"00",	-- Hex Addr	5391	21393
x"00",	-- Hex Addr	5392	21394
x"00",	-- Hex Addr	5393	21395
x"00",	-- Hex Addr	5394	21396
x"00",	-- Hex Addr	5395	21397
x"00",	-- Hex Addr	5396	21398
x"00",	-- Hex Addr	5397	21399
x"00",	-- Hex Addr	5398	21400
x"00",	-- Hex Addr	5399	21401
x"00",	-- Hex Addr	539A	21402
x"00",	-- Hex Addr	539B	21403
x"00",	-- Hex Addr	539C	21404
x"00",	-- Hex Addr	539D	21405
x"00",	-- Hex Addr	539E	21406
x"00",	-- Hex Addr	539F	21407
x"00",	-- Hex Addr	53A0	21408
x"00",	-- Hex Addr	53A1	21409
x"00",	-- Hex Addr	53A2	21410
x"00",	-- Hex Addr	53A3	21411
x"00",	-- Hex Addr	53A4	21412
x"00",	-- Hex Addr	53A5	21413
x"00",	-- Hex Addr	53A6	21414
x"00",	-- Hex Addr	53A7	21415
x"00",	-- Hex Addr	53A8	21416
x"00",	-- Hex Addr	53A9	21417
x"00",	-- Hex Addr	53AA	21418
x"00",	-- Hex Addr	53AB	21419
x"00",	-- Hex Addr	53AC	21420
x"00",	-- Hex Addr	53AD	21421
x"00",	-- Hex Addr	53AE	21422
x"00",	-- Hex Addr	53AF	21423
x"00",	-- Hex Addr	53B0	21424
x"00",	-- Hex Addr	53B1	21425
x"00",	-- Hex Addr	53B2	21426
x"00",	-- Hex Addr	53B3	21427
x"00",	-- Hex Addr	53B4	21428
x"00",	-- Hex Addr	53B5	21429
x"00",	-- Hex Addr	53B6	21430
x"00",	-- Hex Addr	53B7	21431
x"00",	-- Hex Addr	53B8	21432
x"00",	-- Hex Addr	53B9	21433
x"00",	-- Hex Addr	53BA	21434
x"00",	-- Hex Addr	53BB	21435
x"00",	-- Hex Addr	53BC	21436
x"00",	-- Hex Addr	53BD	21437
x"00",	-- Hex Addr	53BE	21438
x"00",	-- Hex Addr	53BF	21439
x"00",	-- Hex Addr	53C0	21440
x"00",	-- Hex Addr	53C1	21441
x"00",	-- Hex Addr	53C2	21442
x"00",	-- Hex Addr	53C3	21443
x"00",	-- Hex Addr	53C4	21444
x"00",	-- Hex Addr	53C5	21445
x"00",	-- Hex Addr	53C6	21446
x"00",	-- Hex Addr	53C7	21447
x"00",	-- Hex Addr	53C8	21448
x"00",	-- Hex Addr	53C9	21449
x"00",	-- Hex Addr	53CA	21450
x"00",	-- Hex Addr	53CB	21451
x"00",	-- Hex Addr	53CC	21452
x"00",	-- Hex Addr	53CD	21453
x"00",	-- Hex Addr	53CE	21454
x"00",	-- Hex Addr	53CF	21455
x"00",	-- Hex Addr	53D0	21456
x"00",	-- Hex Addr	53D1	21457
x"00",	-- Hex Addr	53D2	21458
x"00",	-- Hex Addr	53D3	21459
x"00",	-- Hex Addr	53D4	21460
x"00",	-- Hex Addr	53D5	21461
x"00",	-- Hex Addr	53D6	21462
x"00",	-- Hex Addr	53D7	21463
x"00",	-- Hex Addr	53D8	21464
x"00",	-- Hex Addr	53D9	21465
x"00",	-- Hex Addr	53DA	21466
x"00",	-- Hex Addr	53DB	21467
x"00",	-- Hex Addr	53DC	21468
x"00",	-- Hex Addr	53DD	21469
x"00",	-- Hex Addr	53DE	21470
x"00",	-- Hex Addr	53DF	21471
x"00",	-- Hex Addr	53E0	21472
x"00",	-- Hex Addr	53E1	21473
x"00",	-- Hex Addr	53E2	21474
x"00",	-- Hex Addr	53E3	21475
x"00",	-- Hex Addr	53E4	21476
x"00",	-- Hex Addr	53E5	21477
x"00",	-- Hex Addr	53E6	21478
x"00",	-- Hex Addr	53E7	21479
x"00",	-- Hex Addr	53E8	21480
x"00",	-- Hex Addr	53E9	21481
x"00",	-- Hex Addr	53EA	21482
x"00",	-- Hex Addr	53EB	21483
x"00",	-- Hex Addr	53EC	21484
x"00",	-- Hex Addr	53ED	21485
x"00",	-- Hex Addr	53EE	21486
x"00",	-- Hex Addr	53EF	21487
x"00",	-- Hex Addr	53F0	21488
x"00",	-- Hex Addr	53F1	21489
x"00",	-- Hex Addr	53F2	21490
x"00",	-- Hex Addr	53F3	21491
x"00",	-- Hex Addr	53F4	21492
x"00",	-- Hex Addr	53F5	21493
x"00",	-- Hex Addr	53F6	21494
x"00",	-- Hex Addr	53F7	21495
x"00",	-- Hex Addr	53F8	21496
x"00",	-- Hex Addr	53F9	21497
x"00",	-- Hex Addr	53FA	21498
x"00",	-- Hex Addr	53FB	21499
x"00",	-- Hex Addr	53FC	21500
x"00",	-- Hex Addr	53FD	21501
x"00",	-- Hex Addr	53FE	21502
x"00",	-- Hex Addr	53FF	21503
x"00",	-- Hex Addr	5400	21504
x"00",	-- Hex Addr	5401	21505
x"00",	-- Hex Addr	5402	21506
x"00",	-- Hex Addr	5403	21507
x"00",	-- Hex Addr	5404	21508
x"00",	-- Hex Addr	5405	21509
x"00",	-- Hex Addr	5406	21510
x"00",	-- Hex Addr	5407	21511
x"00",	-- Hex Addr	5408	21512
x"00",	-- Hex Addr	5409	21513
x"00",	-- Hex Addr	540A	21514
x"00",	-- Hex Addr	540B	21515
x"00",	-- Hex Addr	540C	21516
x"00",	-- Hex Addr	540D	21517
x"00",	-- Hex Addr	540E	21518
x"00",	-- Hex Addr	540F	21519
x"00",	-- Hex Addr	5410	21520
x"00",	-- Hex Addr	5411	21521
x"00",	-- Hex Addr	5412	21522
x"00",	-- Hex Addr	5413	21523
x"00",	-- Hex Addr	5414	21524
x"00",	-- Hex Addr	5415	21525
x"00",	-- Hex Addr	5416	21526
x"00",	-- Hex Addr	5417	21527
x"00",	-- Hex Addr	5418	21528
x"00",	-- Hex Addr	5419	21529
x"00",	-- Hex Addr	541A	21530
x"00",	-- Hex Addr	541B	21531
x"00",	-- Hex Addr	541C	21532
x"00",	-- Hex Addr	541D	21533
x"00",	-- Hex Addr	541E	21534
x"00",	-- Hex Addr	541F	21535
x"00",	-- Hex Addr	5420	21536
x"00",	-- Hex Addr	5421	21537
x"00",	-- Hex Addr	5422	21538
x"00",	-- Hex Addr	5423	21539
x"00",	-- Hex Addr	5424	21540
x"00",	-- Hex Addr	5425	21541
x"00",	-- Hex Addr	5426	21542
x"00",	-- Hex Addr	5427	21543
x"00",	-- Hex Addr	5428	21544
x"00",	-- Hex Addr	5429	21545
x"00",	-- Hex Addr	542A	21546
x"00",	-- Hex Addr	542B	21547
x"00",	-- Hex Addr	542C	21548
x"00",	-- Hex Addr	542D	21549
x"00",	-- Hex Addr	542E	21550
x"00",	-- Hex Addr	542F	21551
x"00",	-- Hex Addr	5430	21552
x"00",	-- Hex Addr	5431	21553
x"00",	-- Hex Addr	5432	21554
x"00",	-- Hex Addr	5433	21555
x"00",	-- Hex Addr	5434	21556
x"00",	-- Hex Addr	5435	21557
x"00",	-- Hex Addr	5436	21558
x"00",	-- Hex Addr	5437	21559
x"00",	-- Hex Addr	5438	21560
x"00",	-- Hex Addr	5439	21561
x"00",	-- Hex Addr	543A	21562
x"00",	-- Hex Addr	543B	21563
x"00",	-- Hex Addr	543C	21564
x"00",	-- Hex Addr	543D	21565
x"00",	-- Hex Addr	543E	21566
x"00",	-- Hex Addr	543F	21567
x"00",	-- Hex Addr	5440	21568
x"00",	-- Hex Addr	5441	21569
x"00",	-- Hex Addr	5442	21570
x"00",	-- Hex Addr	5443	21571
x"00",	-- Hex Addr	5444	21572
x"00",	-- Hex Addr	5445	21573
x"00",	-- Hex Addr	5446	21574
x"00",	-- Hex Addr	5447	21575
x"00",	-- Hex Addr	5448	21576
x"00",	-- Hex Addr	5449	21577
x"00",	-- Hex Addr	544A	21578
x"00",	-- Hex Addr	544B	21579
x"00",	-- Hex Addr	544C	21580
x"00",	-- Hex Addr	544D	21581
x"00",	-- Hex Addr	544E	21582
x"00",	-- Hex Addr	544F	21583
x"00",	-- Hex Addr	5450	21584
x"00",	-- Hex Addr	5451	21585
x"00",	-- Hex Addr	5452	21586
x"00",	-- Hex Addr	5453	21587
x"00",	-- Hex Addr	5454	21588
x"00",	-- Hex Addr	5455	21589
x"00",	-- Hex Addr	5456	21590
x"00",	-- Hex Addr	5457	21591
x"00",	-- Hex Addr	5458	21592
x"00",	-- Hex Addr	5459	21593
x"00",	-- Hex Addr	545A	21594
x"00",	-- Hex Addr	545B	21595
x"00",	-- Hex Addr	545C	21596
x"00",	-- Hex Addr	545D	21597
x"00",	-- Hex Addr	545E	21598
x"00",	-- Hex Addr	545F	21599
x"00",	-- Hex Addr	5460	21600
x"00",	-- Hex Addr	5461	21601
x"00",	-- Hex Addr	5462	21602
x"00",	-- Hex Addr	5463	21603
x"00",	-- Hex Addr	5464	21604
x"00",	-- Hex Addr	5465	21605
x"00",	-- Hex Addr	5466	21606
x"00",	-- Hex Addr	5467	21607
x"00",	-- Hex Addr	5468	21608
x"00",	-- Hex Addr	5469	21609
x"00",	-- Hex Addr	546A	21610
x"00",	-- Hex Addr	546B	21611
x"00",	-- Hex Addr	546C	21612
x"00",	-- Hex Addr	546D	21613
x"00",	-- Hex Addr	546E	21614
x"00",	-- Hex Addr	546F	21615
x"00",	-- Hex Addr	5470	21616
x"00",	-- Hex Addr	5471	21617
x"00",	-- Hex Addr	5472	21618
x"00",	-- Hex Addr	5473	21619
x"00",	-- Hex Addr	5474	21620
x"00",	-- Hex Addr	5475	21621
x"00",	-- Hex Addr	5476	21622
x"00",	-- Hex Addr	5477	21623
x"00",	-- Hex Addr	5478	21624
x"00",	-- Hex Addr	5479	21625
x"00",	-- Hex Addr	547A	21626
x"00",	-- Hex Addr	547B	21627
x"00",	-- Hex Addr	547C	21628
x"00",	-- Hex Addr	547D	21629
x"00",	-- Hex Addr	547E	21630
x"00",	-- Hex Addr	547F	21631
x"00",	-- Hex Addr	5480	21632
x"00",	-- Hex Addr	5481	21633
x"00",	-- Hex Addr	5482	21634
x"00",	-- Hex Addr	5483	21635
x"00",	-- Hex Addr	5484	21636
x"00",	-- Hex Addr	5485	21637
x"00",	-- Hex Addr	5486	21638
x"00",	-- Hex Addr	5487	21639
x"00",	-- Hex Addr	5488	21640
x"00",	-- Hex Addr	5489	21641
x"00",	-- Hex Addr	548A	21642
x"00",	-- Hex Addr	548B	21643
x"00",	-- Hex Addr	548C	21644
x"00",	-- Hex Addr	548D	21645
x"00",	-- Hex Addr	548E	21646
x"00",	-- Hex Addr	548F	21647
x"00",	-- Hex Addr	5490	21648
x"00",	-- Hex Addr	5491	21649
x"00",	-- Hex Addr	5492	21650
x"00",	-- Hex Addr	5493	21651
x"00",	-- Hex Addr	5494	21652
x"00",	-- Hex Addr	5495	21653
x"00",	-- Hex Addr	5496	21654
x"00",	-- Hex Addr	5497	21655
x"00",	-- Hex Addr	5498	21656
x"00",	-- Hex Addr	5499	21657
x"00",	-- Hex Addr	549A	21658
x"00",	-- Hex Addr	549B	21659
x"00",	-- Hex Addr	549C	21660
x"00",	-- Hex Addr	549D	21661
x"00",	-- Hex Addr	549E	21662
x"00",	-- Hex Addr	549F	21663
x"00",	-- Hex Addr	54A0	21664
x"00",	-- Hex Addr	54A1	21665
x"00",	-- Hex Addr	54A2	21666
x"00",	-- Hex Addr	54A3	21667
x"00",	-- Hex Addr	54A4	21668
x"00",	-- Hex Addr	54A5	21669
x"00",	-- Hex Addr	54A6	21670
x"00",	-- Hex Addr	54A7	21671
x"00",	-- Hex Addr	54A8	21672
x"00",	-- Hex Addr	54A9	21673
x"00",	-- Hex Addr	54AA	21674
x"00",	-- Hex Addr	54AB	21675
x"00",	-- Hex Addr	54AC	21676
x"00",	-- Hex Addr	54AD	21677
x"00",	-- Hex Addr	54AE	21678
x"00",	-- Hex Addr	54AF	21679
x"00",	-- Hex Addr	54B0	21680
x"00",	-- Hex Addr	54B1	21681
x"00",	-- Hex Addr	54B2	21682
x"00",	-- Hex Addr	54B3	21683
x"00",	-- Hex Addr	54B4	21684
x"00",	-- Hex Addr	54B5	21685
x"00",	-- Hex Addr	54B6	21686
x"00",	-- Hex Addr	54B7	21687
x"00",	-- Hex Addr	54B8	21688
x"00",	-- Hex Addr	54B9	21689
x"00",	-- Hex Addr	54BA	21690
x"00",	-- Hex Addr	54BB	21691
x"00",	-- Hex Addr	54BC	21692
x"00",	-- Hex Addr	54BD	21693
x"00",	-- Hex Addr	54BE	21694
x"00",	-- Hex Addr	54BF	21695
x"00",	-- Hex Addr	54C0	21696
x"00",	-- Hex Addr	54C1	21697
x"00",	-- Hex Addr	54C2	21698
x"00",	-- Hex Addr	54C3	21699
x"00",	-- Hex Addr	54C4	21700
x"00",	-- Hex Addr	54C5	21701
x"00",	-- Hex Addr	54C6	21702
x"00",	-- Hex Addr	54C7	21703
x"00",	-- Hex Addr	54C8	21704
x"00",	-- Hex Addr	54C9	21705
x"00",	-- Hex Addr	54CA	21706
x"00",	-- Hex Addr	54CB	21707
x"00",	-- Hex Addr	54CC	21708
x"00",	-- Hex Addr	54CD	21709
x"00",	-- Hex Addr	54CE	21710
x"00",	-- Hex Addr	54CF	21711
x"00",	-- Hex Addr	54D0	21712
x"00",	-- Hex Addr	54D1	21713
x"00",	-- Hex Addr	54D2	21714
x"00",	-- Hex Addr	54D3	21715
x"00",	-- Hex Addr	54D4	21716
x"00",	-- Hex Addr	54D5	21717
x"00",	-- Hex Addr	54D6	21718
x"00",	-- Hex Addr	54D7	21719
x"00",	-- Hex Addr	54D8	21720
x"00",	-- Hex Addr	54D9	21721
x"00",	-- Hex Addr	54DA	21722
x"00",	-- Hex Addr	54DB	21723
x"00",	-- Hex Addr	54DC	21724
x"00",	-- Hex Addr	54DD	21725
x"00",	-- Hex Addr	54DE	21726
x"00",	-- Hex Addr	54DF	21727
x"00",	-- Hex Addr	54E0	21728
x"00",	-- Hex Addr	54E1	21729
x"00",	-- Hex Addr	54E2	21730
x"00",	-- Hex Addr	54E3	21731
x"00",	-- Hex Addr	54E4	21732
x"00",	-- Hex Addr	54E5	21733
x"00",	-- Hex Addr	54E6	21734
x"00",	-- Hex Addr	54E7	21735
x"00",	-- Hex Addr	54E8	21736
x"00",	-- Hex Addr	54E9	21737
x"00",	-- Hex Addr	54EA	21738
x"00",	-- Hex Addr	54EB	21739
x"00",	-- Hex Addr	54EC	21740
x"00",	-- Hex Addr	54ED	21741
x"00",	-- Hex Addr	54EE	21742
x"00",	-- Hex Addr	54EF	21743
x"00",	-- Hex Addr	54F0	21744
x"00",	-- Hex Addr	54F1	21745
x"00",	-- Hex Addr	54F2	21746
x"00",	-- Hex Addr	54F3	21747
x"00",	-- Hex Addr	54F4	21748
x"00",	-- Hex Addr	54F5	21749
x"00",	-- Hex Addr	54F6	21750
x"00",	-- Hex Addr	54F7	21751
x"00",	-- Hex Addr	54F8	21752
x"00",	-- Hex Addr	54F9	21753
x"00",	-- Hex Addr	54FA	21754
x"00",	-- Hex Addr	54FB	21755
x"00",	-- Hex Addr	54FC	21756
x"00",	-- Hex Addr	54FD	21757
x"00",	-- Hex Addr	54FE	21758
x"00",	-- Hex Addr	54FF	21759
x"00",	-- Hex Addr	5500	21760
x"00",	-- Hex Addr	5501	21761
x"00",	-- Hex Addr	5502	21762
x"00",	-- Hex Addr	5503	21763
x"00",	-- Hex Addr	5504	21764
x"00",	-- Hex Addr	5505	21765
x"00",	-- Hex Addr	5506	21766
x"00",	-- Hex Addr	5507	21767
x"00",	-- Hex Addr	5508	21768
x"00",	-- Hex Addr	5509	21769
x"00",	-- Hex Addr	550A	21770
x"00",	-- Hex Addr	550B	21771
x"00",	-- Hex Addr	550C	21772
x"00",	-- Hex Addr	550D	21773
x"00",	-- Hex Addr	550E	21774
x"00",	-- Hex Addr	550F	21775
x"00",	-- Hex Addr	5510	21776
x"00",	-- Hex Addr	5511	21777
x"00",	-- Hex Addr	5512	21778
x"00",	-- Hex Addr	5513	21779
x"00",	-- Hex Addr	5514	21780
x"00",	-- Hex Addr	5515	21781
x"00",	-- Hex Addr	5516	21782
x"00",	-- Hex Addr	5517	21783
x"00",	-- Hex Addr	5518	21784
x"00",	-- Hex Addr	5519	21785
x"00",	-- Hex Addr	551A	21786
x"00",	-- Hex Addr	551B	21787
x"00",	-- Hex Addr	551C	21788
x"00",	-- Hex Addr	551D	21789
x"00",	-- Hex Addr	551E	21790
x"00",	-- Hex Addr	551F	21791
x"00",	-- Hex Addr	5520	21792
x"00",	-- Hex Addr	5521	21793
x"00",	-- Hex Addr	5522	21794
x"00",	-- Hex Addr	5523	21795
x"00",	-- Hex Addr	5524	21796
x"00",	-- Hex Addr	5525	21797
x"00",	-- Hex Addr	5526	21798
x"00",	-- Hex Addr	5527	21799
x"00",	-- Hex Addr	5528	21800
x"00",	-- Hex Addr	5529	21801
x"00",	-- Hex Addr	552A	21802
x"00",	-- Hex Addr	552B	21803
x"00",	-- Hex Addr	552C	21804
x"00",	-- Hex Addr	552D	21805
x"00",	-- Hex Addr	552E	21806
x"00",	-- Hex Addr	552F	21807
x"00",	-- Hex Addr	5530	21808
x"00",	-- Hex Addr	5531	21809
x"00",	-- Hex Addr	5532	21810
x"00",	-- Hex Addr	5533	21811
x"00",	-- Hex Addr	5534	21812
x"00",	-- Hex Addr	5535	21813
x"00",	-- Hex Addr	5536	21814
x"00",	-- Hex Addr	5537	21815
x"00",	-- Hex Addr	5538	21816
x"00",	-- Hex Addr	5539	21817
x"00",	-- Hex Addr	553A	21818
x"00",	-- Hex Addr	553B	21819
x"00",	-- Hex Addr	553C	21820
x"00",	-- Hex Addr	553D	21821
x"00",	-- Hex Addr	553E	21822
x"00",	-- Hex Addr	553F	21823
x"00",	-- Hex Addr	5540	21824
x"00",	-- Hex Addr	5541	21825
x"00",	-- Hex Addr	5542	21826
x"00",	-- Hex Addr	5543	21827
x"00",	-- Hex Addr	5544	21828
x"00",	-- Hex Addr	5545	21829
x"00",	-- Hex Addr	5546	21830
x"00",	-- Hex Addr	5547	21831
x"00",	-- Hex Addr	5548	21832
x"00",	-- Hex Addr	5549	21833
x"00",	-- Hex Addr	554A	21834
x"00",	-- Hex Addr	554B	21835
x"00",	-- Hex Addr	554C	21836
x"00",	-- Hex Addr	554D	21837
x"00",	-- Hex Addr	554E	21838
x"00",	-- Hex Addr	554F	21839
x"00",	-- Hex Addr	5550	21840
x"00",	-- Hex Addr	5551	21841
x"00",	-- Hex Addr	5552	21842
x"00",	-- Hex Addr	5553	21843
x"00",	-- Hex Addr	5554	21844
x"00",	-- Hex Addr	5555	21845
x"00",	-- Hex Addr	5556	21846
x"00",	-- Hex Addr	5557	21847
x"00",	-- Hex Addr	5558	21848
x"00",	-- Hex Addr	5559	21849
x"00",	-- Hex Addr	555A	21850
x"00",	-- Hex Addr	555B	21851
x"00",	-- Hex Addr	555C	21852
x"00",	-- Hex Addr	555D	21853
x"00",	-- Hex Addr	555E	21854
x"00",	-- Hex Addr	555F	21855
x"00",	-- Hex Addr	5560	21856
x"00",	-- Hex Addr	5561	21857
x"00",	-- Hex Addr	5562	21858
x"00",	-- Hex Addr	5563	21859
x"00",	-- Hex Addr	5564	21860
x"00",	-- Hex Addr	5565	21861
x"00",	-- Hex Addr	5566	21862
x"00",	-- Hex Addr	5567	21863
x"00",	-- Hex Addr	5568	21864
x"00",	-- Hex Addr	5569	21865
x"00",	-- Hex Addr	556A	21866
x"00",	-- Hex Addr	556B	21867
x"00",	-- Hex Addr	556C	21868
x"00",	-- Hex Addr	556D	21869
x"00",	-- Hex Addr	556E	21870
x"00",	-- Hex Addr	556F	21871
x"00",	-- Hex Addr	5570	21872
x"00",	-- Hex Addr	5571	21873
x"00",	-- Hex Addr	5572	21874
x"00",	-- Hex Addr	5573	21875
x"00",	-- Hex Addr	5574	21876
x"00",	-- Hex Addr	5575	21877
x"00",	-- Hex Addr	5576	21878
x"00",	-- Hex Addr	5577	21879
x"00",	-- Hex Addr	5578	21880
x"00",	-- Hex Addr	5579	21881
x"00",	-- Hex Addr	557A	21882
x"00",	-- Hex Addr	557B	21883
x"00",	-- Hex Addr	557C	21884
x"00",	-- Hex Addr	557D	21885
x"00",	-- Hex Addr	557E	21886
x"00",	-- Hex Addr	557F	21887
x"00",	-- Hex Addr	5580	21888
x"00",	-- Hex Addr	5581	21889
x"00",	-- Hex Addr	5582	21890
x"00",	-- Hex Addr	5583	21891
x"00",	-- Hex Addr	5584	21892
x"00",	-- Hex Addr	5585	21893
x"00",	-- Hex Addr	5586	21894
x"00",	-- Hex Addr	5587	21895
x"00",	-- Hex Addr	5588	21896
x"00",	-- Hex Addr	5589	21897
x"00",	-- Hex Addr	558A	21898
x"00",	-- Hex Addr	558B	21899
x"00",	-- Hex Addr	558C	21900
x"00",	-- Hex Addr	558D	21901
x"00",	-- Hex Addr	558E	21902
x"00",	-- Hex Addr	558F	21903
x"00",	-- Hex Addr	5590	21904
x"00",	-- Hex Addr	5591	21905
x"00",	-- Hex Addr	5592	21906
x"00",	-- Hex Addr	5593	21907
x"00",	-- Hex Addr	5594	21908
x"00",	-- Hex Addr	5595	21909
x"00",	-- Hex Addr	5596	21910
x"00",	-- Hex Addr	5597	21911
x"00",	-- Hex Addr	5598	21912
x"00",	-- Hex Addr	5599	21913
x"00",	-- Hex Addr	559A	21914
x"00",	-- Hex Addr	559B	21915
x"00",	-- Hex Addr	559C	21916
x"00",	-- Hex Addr	559D	21917
x"00",	-- Hex Addr	559E	21918
x"00",	-- Hex Addr	559F	21919
x"00",	-- Hex Addr	55A0	21920
x"00",	-- Hex Addr	55A1	21921
x"00",	-- Hex Addr	55A2	21922
x"00",	-- Hex Addr	55A3	21923
x"00",	-- Hex Addr	55A4	21924
x"00",	-- Hex Addr	55A5	21925
x"00",	-- Hex Addr	55A6	21926
x"00",	-- Hex Addr	55A7	21927
x"00",	-- Hex Addr	55A8	21928
x"00",	-- Hex Addr	55A9	21929
x"00",	-- Hex Addr	55AA	21930
x"00",	-- Hex Addr	55AB	21931
x"00",	-- Hex Addr	55AC	21932
x"00",	-- Hex Addr	55AD	21933
x"00",	-- Hex Addr	55AE	21934
x"00",	-- Hex Addr	55AF	21935
x"00",	-- Hex Addr	55B0	21936
x"00",	-- Hex Addr	55B1	21937
x"00",	-- Hex Addr	55B2	21938
x"00",	-- Hex Addr	55B3	21939
x"00",	-- Hex Addr	55B4	21940
x"00",	-- Hex Addr	55B5	21941
x"00",	-- Hex Addr	55B6	21942
x"00",	-- Hex Addr	55B7	21943
x"00",	-- Hex Addr	55B8	21944
x"00",	-- Hex Addr	55B9	21945
x"00",	-- Hex Addr	55BA	21946
x"00",	-- Hex Addr	55BB	21947
x"00",	-- Hex Addr	55BC	21948
x"00",	-- Hex Addr	55BD	21949
x"00",	-- Hex Addr	55BE	21950
x"00",	-- Hex Addr	55BF	21951
x"00",	-- Hex Addr	55C0	21952
x"00",	-- Hex Addr	55C1	21953
x"00",	-- Hex Addr	55C2	21954
x"00",	-- Hex Addr	55C3	21955
x"00",	-- Hex Addr	55C4	21956
x"00",	-- Hex Addr	55C5	21957
x"00",	-- Hex Addr	55C6	21958
x"00",	-- Hex Addr	55C7	21959
x"00",	-- Hex Addr	55C8	21960
x"00",	-- Hex Addr	55C9	21961
x"00",	-- Hex Addr	55CA	21962
x"00",	-- Hex Addr	55CB	21963
x"00",	-- Hex Addr	55CC	21964
x"00",	-- Hex Addr	55CD	21965
x"00",	-- Hex Addr	55CE	21966
x"00",	-- Hex Addr	55CF	21967
x"00",	-- Hex Addr	55D0	21968
x"00",	-- Hex Addr	55D1	21969
x"00",	-- Hex Addr	55D2	21970
x"00",	-- Hex Addr	55D3	21971
x"00",	-- Hex Addr	55D4	21972
x"00",	-- Hex Addr	55D5	21973
x"00",	-- Hex Addr	55D6	21974
x"00",	-- Hex Addr	55D7	21975
x"00",	-- Hex Addr	55D8	21976
x"00",	-- Hex Addr	55D9	21977
x"00",	-- Hex Addr	55DA	21978
x"00",	-- Hex Addr	55DB	21979
x"00",	-- Hex Addr	55DC	21980
x"00",	-- Hex Addr	55DD	21981
x"00",	-- Hex Addr	55DE	21982
x"00",	-- Hex Addr	55DF	21983
x"00",	-- Hex Addr	55E0	21984
x"00",	-- Hex Addr	55E1	21985
x"00",	-- Hex Addr	55E2	21986
x"00",	-- Hex Addr	55E3	21987
x"00",	-- Hex Addr	55E4	21988
x"00",	-- Hex Addr	55E5	21989
x"00",	-- Hex Addr	55E6	21990
x"00",	-- Hex Addr	55E7	21991
x"00",	-- Hex Addr	55E8	21992
x"00",	-- Hex Addr	55E9	21993
x"00",	-- Hex Addr	55EA	21994
x"00",	-- Hex Addr	55EB	21995
x"00",	-- Hex Addr	55EC	21996
x"00",	-- Hex Addr	55ED	21997
x"00",	-- Hex Addr	55EE	21998
x"00",	-- Hex Addr	55EF	21999
x"00",	-- Hex Addr	55F0	22000
x"00",	-- Hex Addr	55F1	22001
x"00",	-- Hex Addr	55F2	22002
x"00",	-- Hex Addr	55F3	22003
x"00",	-- Hex Addr	55F4	22004
x"00",	-- Hex Addr	55F5	22005
x"00",	-- Hex Addr	55F6	22006
x"00",	-- Hex Addr	55F7	22007
x"00",	-- Hex Addr	55F8	22008
x"00",	-- Hex Addr	55F9	22009
x"00",	-- Hex Addr	55FA	22010
x"00",	-- Hex Addr	55FB	22011
x"00",	-- Hex Addr	55FC	22012
x"00",	-- Hex Addr	55FD	22013
x"00",	-- Hex Addr	55FE	22014
x"00",	-- Hex Addr	55FF	22015
x"00",	-- Hex Addr	5600	22016
x"00",	-- Hex Addr	5601	22017
x"00",	-- Hex Addr	5602	22018
x"00",	-- Hex Addr	5603	22019
x"00",	-- Hex Addr	5604	22020
x"00",	-- Hex Addr	5605	22021
x"00",	-- Hex Addr	5606	22022
x"00",	-- Hex Addr	5607	22023
x"00",	-- Hex Addr	5608	22024
x"00",	-- Hex Addr	5609	22025
x"00",	-- Hex Addr	560A	22026
x"00",	-- Hex Addr	560B	22027
x"00",	-- Hex Addr	560C	22028
x"00",	-- Hex Addr	560D	22029
x"00",	-- Hex Addr	560E	22030
x"00",	-- Hex Addr	560F	22031
x"00",	-- Hex Addr	5610	22032
x"00",	-- Hex Addr	5611	22033
x"00",	-- Hex Addr	5612	22034
x"00",	-- Hex Addr	5613	22035
x"00",	-- Hex Addr	5614	22036
x"00",	-- Hex Addr	5615	22037
x"00",	-- Hex Addr	5616	22038
x"00",	-- Hex Addr	5617	22039
x"00",	-- Hex Addr	5618	22040
x"00",	-- Hex Addr	5619	22041
x"00",	-- Hex Addr	561A	22042
x"00",	-- Hex Addr	561B	22043
x"00",	-- Hex Addr	561C	22044
x"00",	-- Hex Addr	561D	22045
x"00",	-- Hex Addr	561E	22046
x"00",	-- Hex Addr	561F	22047
x"00",	-- Hex Addr	5620	22048
x"00",	-- Hex Addr	5621	22049
x"00",	-- Hex Addr	5622	22050
x"00",	-- Hex Addr	5623	22051
x"00",	-- Hex Addr	5624	22052
x"00",	-- Hex Addr	5625	22053
x"00",	-- Hex Addr	5626	22054
x"00",	-- Hex Addr	5627	22055
x"00",	-- Hex Addr	5628	22056
x"00",	-- Hex Addr	5629	22057
x"00",	-- Hex Addr	562A	22058
x"00",	-- Hex Addr	562B	22059
x"00",	-- Hex Addr	562C	22060
x"00",	-- Hex Addr	562D	22061
x"00",	-- Hex Addr	562E	22062
x"00",	-- Hex Addr	562F	22063
x"00",	-- Hex Addr	5630	22064
x"00",	-- Hex Addr	5631	22065
x"00",	-- Hex Addr	5632	22066
x"00",	-- Hex Addr	5633	22067
x"00",	-- Hex Addr	5634	22068
x"00",	-- Hex Addr	5635	22069
x"00",	-- Hex Addr	5636	22070
x"00",	-- Hex Addr	5637	22071
x"00",	-- Hex Addr	5638	22072
x"00",	-- Hex Addr	5639	22073
x"00",	-- Hex Addr	563A	22074
x"00",	-- Hex Addr	563B	22075
x"00",	-- Hex Addr	563C	22076
x"00",	-- Hex Addr	563D	22077
x"00",	-- Hex Addr	563E	22078
x"00",	-- Hex Addr	563F	22079
x"00",	-- Hex Addr	5640	22080
x"00",	-- Hex Addr	5641	22081
x"00",	-- Hex Addr	5642	22082
x"00",	-- Hex Addr	5643	22083
x"00",	-- Hex Addr	5644	22084
x"00",	-- Hex Addr	5645	22085
x"00",	-- Hex Addr	5646	22086
x"00",	-- Hex Addr	5647	22087
x"00",	-- Hex Addr	5648	22088
x"00",	-- Hex Addr	5649	22089
x"00",	-- Hex Addr	564A	22090
x"00",	-- Hex Addr	564B	22091
x"00",	-- Hex Addr	564C	22092
x"00",	-- Hex Addr	564D	22093
x"00",	-- Hex Addr	564E	22094
x"00",	-- Hex Addr	564F	22095
x"00",	-- Hex Addr	5650	22096
x"00",	-- Hex Addr	5651	22097
x"00",	-- Hex Addr	5652	22098
x"00",	-- Hex Addr	5653	22099
x"00",	-- Hex Addr	5654	22100
x"00",	-- Hex Addr	5655	22101
x"00",	-- Hex Addr	5656	22102
x"00",	-- Hex Addr	5657	22103
x"00",	-- Hex Addr	5658	22104
x"00",	-- Hex Addr	5659	22105
x"00",	-- Hex Addr	565A	22106
x"00",	-- Hex Addr	565B	22107
x"00",	-- Hex Addr	565C	22108
x"00",	-- Hex Addr	565D	22109
x"00",	-- Hex Addr	565E	22110
x"00",	-- Hex Addr	565F	22111
x"00",	-- Hex Addr	5660	22112
x"00",	-- Hex Addr	5661	22113
x"00",	-- Hex Addr	5662	22114
x"00",	-- Hex Addr	5663	22115
x"00",	-- Hex Addr	5664	22116
x"00",	-- Hex Addr	5665	22117
x"00",	-- Hex Addr	5666	22118
x"00",	-- Hex Addr	5667	22119
x"00",	-- Hex Addr	5668	22120
x"00",	-- Hex Addr	5669	22121
x"00",	-- Hex Addr	566A	22122
x"00",	-- Hex Addr	566B	22123
x"00",	-- Hex Addr	566C	22124
x"00",	-- Hex Addr	566D	22125
x"00",	-- Hex Addr	566E	22126
x"00",	-- Hex Addr	566F	22127
x"00",	-- Hex Addr	5670	22128
x"00",	-- Hex Addr	5671	22129
x"00",	-- Hex Addr	5672	22130
x"00",	-- Hex Addr	5673	22131
x"00",	-- Hex Addr	5674	22132
x"00",	-- Hex Addr	5675	22133
x"00",	-- Hex Addr	5676	22134
x"00",	-- Hex Addr	5677	22135
x"00",	-- Hex Addr	5678	22136
x"00",	-- Hex Addr	5679	22137
x"00",	-- Hex Addr	567A	22138
x"00",	-- Hex Addr	567B	22139
x"00",	-- Hex Addr	567C	22140
x"00",	-- Hex Addr	567D	22141
x"00",	-- Hex Addr	567E	22142
x"00",	-- Hex Addr	567F	22143
x"00",	-- Hex Addr	5680	22144
x"00",	-- Hex Addr	5681	22145
x"00",	-- Hex Addr	5682	22146
x"00",	-- Hex Addr	5683	22147
x"00",	-- Hex Addr	5684	22148
x"00",	-- Hex Addr	5685	22149
x"00",	-- Hex Addr	5686	22150
x"00",	-- Hex Addr	5687	22151
x"00",	-- Hex Addr	5688	22152
x"00",	-- Hex Addr	5689	22153
x"00",	-- Hex Addr	568A	22154
x"00",	-- Hex Addr	568B	22155
x"00",	-- Hex Addr	568C	22156
x"00",	-- Hex Addr	568D	22157
x"00",	-- Hex Addr	568E	22158
x"00",	-- Hex Addr	568F	22159
x"00",	-- Hex Addr	5690	22160
x"00",	-- Hex Addr	5691	22161
x"00",	-- Hex Addr	5692	22162
x"00",	-- Hex Addr	5693	22163
x"00",	-- Hex Addr	5694	22164
x"00",	-- Hex Addr	5695	22165
x"00",	-- Hex Addr	5696	22166
x"00",	-- Hex Addr	5697	22167
x"00",	-- Hex Addr	5698	22168
x"00",	-- Hex Addr	5699	22169
x"00",	-- Hex Addr	569A	22170
x"00",	-- Hex Addr	569B	22171
x"00",	-- Hex Addr	569C	22172
x"00",	-- Hex Addr	569D	22173
x"00",	-- Hex Addr	569E	22174
x"00",	-- Hex Addr	569F	22175
x"00",	-- Hex Addr	56A0	22176
x"00",	-- Hex Addr	56A1	22177
x"00",	-- Hex Addr	56A2	22178
x"00",	-- Hex Addr	56A3	22179
x"00",	-- Hex Addr	56A4	22180
x"00",	-- Hex Addr	56A5	22181
x"00",	-- Hex Addr	56A6	22182
x"00",	-- Hex Addr	56A7	22183
x"00",	-- Hex Addr	56A8	22184
x"00",	-- Hex Addr	56A9	22185
x"00",	-- Hex Addr	56AA	22186
x"00",	-- Hex Addr	56AB	22187
x"00",	-- Hex Addr	56AC	22188
x"00",	-- Hex Addr	56AD	22189
x"00",	-- Hex Addr	56AE	22190
x"00",	-- Hex Addr	56AF	22191
x"00",	-- Hex Addr	56B0	22192
x"00",	-- Hex Addr	56B1	22193
x"00",	-- Hex Addr	56B2	22194
x"00",	-- Hex Addr	56B3	22195
x"00",	-- Hex Addr	56B4	22196
x"00",	-- Hex Addr	56B5	22197
x"00",	-- Hex Addr	56B6	22198
x"00",	-- Hex Addr	56B7	22199
x"00",	-- Hex Addr	56B8	22200
x"00",	-- Hex Addr	56B9	22201
x"00",	-- Hex Addr	56BA	22202
x"00",	-- Hex Addr	56BB	22203
x"00",	-- Hex Addr	56BC	22204
x"00",	-- Hex Addr	56BD	22205
x"00",	-- Hex Addr	56BE	22206
x"00",	-- Hex Addr	56BF	22207
x"00",	-- Hex Addr	56C0	22208
x"00",	-- Hex Addr	56C1	22209
x"00",	-- Hex Addr	56C2	22210
x"00",	-- Hex Addr	56C3	22211
x"00",	-- Hex Addr	56C4	22212
x"00",	-- Hex Addr	56C5	22213
x"00",	-- Hex Addr	56C6	22214
x"00",	-- Hex Addr	56C7	22215
x"00",	-- Hex Addr	56C8	22216
x"00",	-- Hex Addr	56C9	22217
x"00",	-- Hex Addr	56CA	22218
x"00",	-- Hex Addr	56CB	22219
x"00",	-- Hex Addr	56CC	22220
x"00",	-- Hex Addr	56CD	22221
x"00",	-- Hex Addr	56CE	22222
x"00",	-- Hex Addr	56CF	22223
x"00",	-- Hex Addr	56D0	22224
x"00",	-- Hex Addr	56D1	22225
x"00",	-- Hex Addr	56D2	22226
x"00",	-- Hex Addr	56D3	22227
x"00",	-- Hex Addr	56D4	22228
x"00",	-- Hex Addr	56D5	22229
x"00",	-- Hex Addr	56D6	22230
x"00",	-- Hex Addr	56D7	22231
x"00",	-- Hex Addr	56D8	22232
x"00",	-- Hex Addr	56D9	22233
x"00",	-- Hex Addr	56DA	22234
x"00",	-- Hex Addr	56DB	22235
x"00",	-- Hex Addr	56DC	22236
x"00",	-- Hex Addr	56DD	22237
x"00",	-- Hex Addr	56DE	22238
x"00",	-- Hex Addr	56DF	22239
x"00",	-- Hex Addr	56E0	22240
x"00",	-- Hex Addr	56E1	22241
x"00",	-- Hex Addr	56E2	22242
x"00",	-- Hex Addr	56E3	22243
x"00",	-- Hex Addr	56E4	22244
x"00",	-- Hex Addr	56E5	22245
x"00",	-- Hex Addr	56E6	22246
x"00",	-- Hex Addr	56E7	22247
x"00",	-- Hex Addr	56E8	22248
x"00",	-- Hex Addr	56E9	22249
x"00",	-- Hex Addr	56EA	22250
x"00",	-- Hex Addr	56EB	22251
x"00",	-- Hex Addr	56EC	22252
x"00",	-- Hex Addr	56ED	22253
x"00",	-- Hex Addr	56EE	22254
x"00",	-- Hex Addr	56EF	22255
x"00",	-- Hex Addr	56F0	22256
x"00",	-- Hex Addr	56F1	22257
x"00",	-- Hex Addr	56F2	22258
x"00",	-- Hex Addr	56F3	22259
x"00",	-- Hex Addr	56F4	22260
x"00",	-- Hex Addr	56F5	22261
x"00",	-- Hex Addr	56F6	22262
x"00",	-- Hex Addr	56F7	22263
x"00",	-- Hex Addr	56F8	22264
x"00",	-- Hex Addr	56F9	22265
x"00",	-- Hex Addr	56FA	22266
x"00",	-- Hex Addr	56FB	22267
x"00",	-- Hex Addr	56FC	22268
x"00",	-- Hex Addr	56FD	22269
x"00",	-- Hex Addr	56FE	22270
x"00",	-- Hex Addr	56FF	22271
x"00",	-- Hex Addr	5700	22272
x"00",	-- Hex Addr	5701	22273
x"00",	-- Hex Addr	5702	22274
x"00",	-- Hex Addr	5703	22275
x"00",	-- Hex Addr	5704	22276
x"00",	-- Hex Addr	5705	22277
x"00",	-- Hex Addr	5706	22278
x"00",	-- Hex Addr	5707	22279
x"00",	-- Hex Addr	5708	22280
x"00",	-- Hex Addr	5709	22281
x"00",	-- Hex Addr	570A	22282
x"00",	-- Hex Addr	570B	22283
x"00",	-- Hex Addr	570C	22284
x"00",	-- Hex Addr	570D	22285
x"00",	-- Hex Addr	570E	22286
x"00",	-- Hex Addr	570F	22287
x"00",	-- Hex Addr	5710	22288
x"00",	-- Hex Addr	5711	22289
x"00",	-- Hex Addr	5712	22290
x"00",	-- Hex Addr	5713	22291
x"00",	-- Hex Addr	5714	22292
x"00",	-- Hex Addr	5715	22293
x"00",	-- Hex Addr	5716	22294
x"00",	-- Hex Addr	5717	22295
x"00",	-- Hex Addr	5718	22296
x"00",	-- Hex Addr	5719	22297
x"00",	-- Hex Addr	571A	22298
x"00",	-- Hex Addr	571B	22299
x"00",	-- Hex Addr	571C	22300
x"00",	-- Hex Addr	571D	22301
x"00",	-- Hex Addr	571E	22302
x"00",	-- Hex Addr	571F	22303
x"00",	-- Hex Addr	5720	22304
x"00",	-- Hex Addr	5721	22305
x"00",	-- Hex Addr	5722	22306
x"00",	-- Hex Addr	5723	22307
x"00",	-- Hex Addr	5724	22308
x"00",	-- Hex Addr	5725	22309
x"00",	-- Hex Addr	5726	22310
x"00",	-- Hex Addr	5727	22311
x"00",	-- Hex Addr	5728	22312
x"00",	-- Hex Addr	5729	22313
x"00",	-- Hex Addr	572A	22314
x"00",	-- Hex Addr	572B	22315
x"00",	-- Hex Addr	572C	22316
x"00",	-- Hex Addr	572D	22317
x"00",	-- Hex Addr	572E	22318
x"00",	-- Hex Addr	572F	22319
x"00",	-- Hex Addr	5730	22320
x"00",	-- Hex Addr	5731	22321
x"00",	-- Hex Addr	5732	22322
x"00",	-- Hex Addr	5733	22323
x"00",	-- Hex Addr	5734	22324
x"00",	-- Hex Addr	5735	22325
x"00",	-- Hex Addr	5736	22326
x"00",	-- Hex Addr	5737	22327
x"00",	-- Hex Addr	5738	22328
x"00",	-- Hex Addr	5739	22329
x"00",	-- Hex Addr	573A	22330
x"00",	-- Hex Addr	573B	22331
x"00",	-- Hex Addr	573C	22332
x"00",	-- Hex Addr	573D	22333
x"00",	-- Hex Addr	573E	22334
x"00",	-- Hex Addr	573F	22335
x"00",	-- Hex Addr	5740	22336
x"00",	-- Hex Addr	5741	22337
x"00",	-- Hex Addr	5742	22338
x"00",	-- Hex Addr	5743	22339
x"00",	-- Hex Addr	5744	22340
x"00",	-- Hex Addr	5745	22341
x"00",	-- Hex Addr	5746	22342
x"00",	-- Hex Addr	5747	22343
x"00",	-- Hex Addr	5748	22344
x"00",	-- Hex Addr	5749	22345
x"00",	-- Hex Addr	574A	22346
x"00",	-- Hex Addr	574B	22347
x"00",	-- Hex Addr	574C	22348
x"00",	-- Hex Addr	574D	22349
x"00",	-- Hex Addr	574E	22350
x"00",	-- Hex Addr	574F	22351
x"00",	-- Hex Addr	5750	22352
x"00",	-- Hex Addr	5751	22353
x"00",	-- Hex Addr	5752	22354
x"00",	-- Hex Addr	5753	22355
x"00",	-- Hex Addr	5754	22356
x"00",	-- Hex Addr	5755	22357
x"00",	-- Hex Addr	5756	22358
x"00",	-- Hex Addr	5757	22359
x"00",	-- Hex Addr	5758	22360
x"00",	-- Hex Addr	5759	22361
x"00",	-- Hex Addr	575A	22362
x"00",	-- Hex Addr	575B	22363
x"00",	-- Hex Addr	575C	22364
x"00",	-- Hex Addr	575D	22365
x"00",	-- Hex Addr	575E	22366
x"00",	-- Hex Addr	575F	22367
x"00",	-- Hex Addr	5760	22368
x"00",	-- Hex Addr	5761	22369
x"00",	-- Hex Addr	5762	22370
x"00",	-- Hex Addr	5763	22371
x"00",	-- Hex Addr	5764	22372
x"00",	-- Hex Addr	5765	22373
x"00",	-- Hex Addr	5766	22374
x"00",	-- Hex Addr	5767	22375
x"00",	-- Hex Addr	5768	22376
x"00",	-- Hex Addr	5769	22377
x"00",	-- Hex Addr	576A	22378
x"00",	-- Hex Addr	576B	22379
x"00",	-- Hex Addr	576C	22380
x"00",	-- Hex Addr	576D	22381
x"00",	-- Hex Addr	576E	22382
x"00",	-- Hex Addr	576F	22383
x"00",	-- Hex Addr	5770	22384
x"00",	-- Hex Addr	5771	22385
x"00",	-- Hex Addr	5772	22386
x"00",	-- Hex Addr	5773	22387
x"00",	-- Hex Addr	5774	22388
x"00",	-- Hex Addr	5775	22389
x"00",	-- Hex Addr	5776	22390
x"00",	-- Hex Addr	5777	22391
x"00",	-- Hex Addr	5778	22392
x"00",	-- Hex Addr	5779	22393
x"00",	-- Hex Addr	577A	22394
x"00",	-- Hex Addr	577B	22395
x"00",	-- Hex Addr	577C	22396
x"00",	-- Hex Addr	577D	22397
x"00",	-- Hex Addr	577E	22398
x"00",	-- Hex Addr	577F	22399
x"00",	-- Hex Addr	5780	22400
x"00",	-- Hex Addr	5781	22401
x"00",	-- Hex Addr	5782	22402
x"00",	-- Hex Addr	5783	22403
x"00",	-- Hex Addr	5784	22404
x"00",	-- Hex Addr	5785	22405
x"00",	-- Hex Addr	5786	22406
x"00",	-- Hex Addr	5787	22407
x"00",	-- Hex Addr	5788	22408
x"00",	-- Hex Addr	5789	22409
x"00",	-- Hex Addr	578A	22410
x"00",	-- Hex Addr	578B	22411
x"00",	-- Hex Addr	578C	22412
x"00",	-- Hex Addr	578D	22413
x"00",	-- Hex Addr	578E	22414
x"00",	-- Hex Addr	578F	22415
x"00",	-- Hex Addr	5790	22416
x"00",	-- Hex Addr	5791	22417
x"00",	-- Hex Addr	5792	22418
x"00",	-- Hex Addr	5793	22419
x"00",	-- Hex Addr	5794	22420
x"00",	-- Hex Addr	5795	22421
x"00",	-- Hex Addr	5796	22422
x"00",	-- Hex Addr	5797	22423
x"00",	-- Hex Addr	5798	22424
x"00",	-- Hex Addr	5799	22425
x"00",	-- Hex Addr	579A	22426
x"00",	-- Hex Addr	579B	22427
x"00",	-- Hex Addr	579C	22428
x"00",	-- Hex Addr	579D	22429
x"00",	-- Hex Addr	579E	22430
x"00",	-- Hex Addr	579F	22431
x"00",	-- Hex Addr	57A0	22432
x"00",	-- Hex Addr	57A1	22433
x"00",	-- Hex Addr	57A2	22434
x"00",	-- Hex Addr	57A3	22435
x"00",	-- Hex Addr	57A4	22436
x"00",	-- Hex Addr	57A5	22437
x"00",	-- Hex Addr	57A6	22438
x"00",	-- Hex Addr	57A7	22439
x"00",	-- Hex Addr	57A8	22440
x"00",	-- Hex Addr	57A9	22441
x"00",	-- Hex Addr	57AA	22442
x"00",	-- Hex Addr	57AB	22443
x"00",	-- Hex Addr	57AC	22444
x"00",	-- Hex Addr	57AD	22445
x"00",	-- Hex Addr	57AE	22446
x"00",	-- Hex Addr	57AF	22447
x"00",	-- Hex Addr	57B0	22448
x"00",	-- Hex Addr	57B1	22449
x"00",	-- Hex Addr	57B2	22450
x"00",	-- Hex Addr	57B3	22451
x"00",	-- Hex Addr	57B4	22452
x"00",	-- Hex Addr	57B5	22453
x"00",	-- Hex Addr	57B6	22454
x"00",	-- Hex Addr	57B7	22455
x"00",	-- Hex Addr	57B8	22456
x"00",	-- Hex Addr	57B9	22457
x"00",	-- Hex Addr	57BA	22458
x"00",	-- Hex Addr	57BB	22459
x"00",	-- Hex Addr	57BC	22460
x"00",	-- Hex Addr	57BD	22461
x"00",	-- Hex Addr	57BE	22462
x"00",	-- Hex Addr	57BF	22463
x"00",	-- Hex Addr	57C0	22464
x"00",	-- Hex Addr	57C1	22465
x"00",	-- Hex Addr	57C2	22466
x"00",	-- Hex Addr	57C3	22467
x"00",	-- Hex Addr	57C4	22468
x"00",	-- Hex Addr	57C5	22469
x"00",	-- Hex Addr	57C6	22470
x"00",	-- Hex Addr	57C7	22471
x"00",	-- Hex Addr	57C8	22472
x"00",	-- Hex Addr	57C9	22473
x"00",	-- Hex Addr	57CA	22474
x"00",	-- Hex Addr	57CB	22475
x"00",	-- Hex Addr	57CC	22476
x"00",	-- Hex Addr	57CD	22477
x"00",	-- Hex Addr	57CE	22478
x"00",	-- Hex Addr	57CF	22479
x"00",	-- Hex Addr	57D0	22480
x"00",	-- Hex Addr	57D1	22481
x"00",	-- Hex Addr	57D2	22482
x"00",	-- Hex Addr	57D3	22483
x"00",	-- Hex Addr	57D4	22484
x"00",	-- Hex Addr	57D5	22485
x"00",	-- Hex Addr	57D6	22486
x"00",	-- Hex Addr	57D7	22487
x"00",	-- Hex Addr	57D8	22488
x"00",	-- Hex Addr	57D9	22489
x"00",	-- Hex Addr	57DA	22490
x"00",	-- Hex Addr	57DB	22491
x"00",	-- Hex Addr	57DC	22492
x"00",	-- Hex Addr	57DD	22493
x"00",	-- Hex Addr	57DE	22494
x"00",	-- Hex Addr	57DF	22495
x"00",	-- Hex Addr	57E0	22496
x"00",	-- Hex Addr	57E1	22497
x"00",	-- Hex Addr	57E2	22498
x"00",	-- Hex Addr	57E3	22499
x"00",	-- Hex Addr	57E4	22500
x"00",	-- Hex Addr	57E5	22501
x"00",	-- Hex Addr	57E6	22502
x"00",	-- Hex Addr	57E7	22503
x"00",	-- Hex Addr	57E8	22504
x"00",	-- Hex Addr	57E9	22505
x"00",	-- Hex Addr	57EA	22506
x"00",	-- Hex Addr	57EB	22507
x"00",	-- Hex Addr	57EC	22508
x"00",	-- Hex Addr	57ED	22509
x"00",	-- Hex Addr	57EE	22510
x"00",	-- Hex Addr	57EF	22511
x"00",	-- Hex Addr	57F0	22512
x"00",	-- Hex Addr	57F1	22513
x"00",	-- Hex Addr	57F2	22514
x"00",	-- Hex Addr	57F3	22515
x"00",	-- Hex Addr	57F4	22516
x"00",	-- Hex Addr	57F5	22517
x"00",	-- Hex Addr	57F6	22518
x"00",	-- Hex Addr	57F7	22519
x"00",	-- Hex Addr	57F8	22520
x"00",	-- Hex Addr	57F9	22521
x"00",	-- Hex Addr	57FA	22522
x"00",	-- Hex Addr	57FB	22523
x"00",	-- Hex Addr	57FC	22524
x"00",	-- Hex Addr	57FD	22525
x"00",	-- Hex Addr	57FE	22526
x"00",	-- Hex Addr	57FF	22527
x"00",	-- Hex Addr	5800	22528
x"00",	-- Hex Addr	5801	22529
x"00",	-- Hex Addr	5802	22530
x"00",	-- Hex Addr	5803	22531
x"00",	-- Hex Addr	5804	22532
x"00",	-- Hex Addr	5805	22533
x"00",	-- Hex Addr	5806	22534
x"00",	-- Hex Addr	5807	22535
x"00",	-- Hex Addr	5808	22536
x"00",	-- Hex Addr	5809	22537
x"00",	-- Hex Addr	580A	22538
x"00",	-- Hex Addr	580B	22539
x"00",	-- Hex Addr	580C	22540
x"00",	-- Hex Addr	580D	22541
x"00",	-- Hex Addr	580E	22542
x"00",	-- Hex Addr	580F	22543
x"00",	-- Hex Addr	5810	22544
x"00",	-- Hex Addr	5811	22545
x"00",	-- Hex Addr	5812	22546
x"00",	-- Hex Addr	5813	22547
x"00",	-- Hex Addr	5814	22548
x"00",	-- Hex Addr	5815	22549
x"00",	-- Hex Addr	5816	22550
x"00",	-- Hex Addr	5817	22551
x"00",	-- Hex Addr	5818	22552
x"00",	-- Hex Addr	5819	22553
x"00",	-- Hex Addr	581A	22554
x"00",	-- Hex Addr	581B	22555
x"00",	-- Hex Addr	581C	22556
x"00",	-- Hex Addr	581D	22557
x"00",	-- Hex Addr	581E	22558
x"00",	-- Hex Addr	581F	22559
x"00",	-- Hex Addr	5820	22560
x"00",	-- Hex Addr	5821	22561
x"00",	-- Hex Addr	5822	22562
x"00",	-- Hex Addr	5823	22563
x"00",	-- Hex Addr	5824	22564
x"00",	-- Hex Addr	5825	22565
x"00",	-- Hex Addr	5826	22566
x"00",	-- Hex Addr	5827	22567
x"00",	-- Hex Addr	5828	22568
x"00",	-- Hex Addr	5829	22569
x"00",	-- Hex Addr	582A	22570
x"00",	-- Hex Addr	582B	22571
x"00",	-- Hex Addr	582C	22572
x"00",	-- Hex Addr	582D	22573
x"00",	-- Hex Addr	582E	22574
x"00",	-- Hex Addr	582F	22575
x"00",	-- Hex Addr	5830	22576
x"00",	-- Hex Addr	5831	22577
x"00",	-- Hex Addr	5832	22578
x"00",	-- Hex Addr	5833	22579
x"00",	-- Hex Addr	5834	22580
x"00",	-- Hex Addr	5835	22581
x"00",	-- Hex Addr	5836	22582
x"00",	-- Hex Addr	5837	22583
x"00",	-- Hex Addr	5838	22584
x"00",	-- Hex Addr	5839	22585
x"00",	-- Hex Addr	583A	22586
x"00",	-- Hex Addr	583B	22587
x"00",	-- Hex Addr	583C	22588
x"00",	-- Hex Addr	583D	22589
x"00",	-- Hex Addr	583E	22590
x"00",	-- Hex Addr	583F	22591
x"00",	-- Hex Addr	5840	22592
x"00",	-- Hex Addr	5841	22593
x"00",	-- Hex Addr	5842	22594
x"00",	-- Hex Addr	5843	22595
x"00",	-- Hex Addr	5844	22596
x"00",	-- Hex Addr	5845	22597
x"00",	-- Hex Addr	5846	22598
x"00",	-- Hex Addr	5847	22599
x"00",	-- Hex Addr	5848	22600
x"00",	-- Hex Addr	5849	22601
x"00",	-- Hex Addr	584A	22602
x"00",	-- Hex Addr	584B	22603
x"00",	-- Hex Addr	584C	22604
x"00",	-- Hex Addr	584D	22605
x"00",	-- Hex Addr	584E	22606
x"00",	-- Hex Addr	584F	22607
x"00",	-- Hex Addr	5850	22608
x"00",	-- Hex Addr	5851	22609
x"00",	-- Hex Addr	5852	22610
x"00",	-- Hex Addr	5853	22611
x"00",	-- Hex Addr	5854	22612
x"00",	-- Hex Addr	5855	22613
x"00",	-- Hex Addr	5856	22614
x"00",	-- Hex Addr	5857	22615
x"00",	-- Hex Addr	5858	22616
x"00",	-- Hex Addr	5859	22617
x"00",	-- Hex Addr	585A	22618
x"00",	-- Hex Addr	585B	22619
x"00",	-- Hex Addr	585C	22620
x"00",	-- Hex Addr	585D	22621
x"00",	-- Hex Addr	585E	22622
x"00",	-- Hex Addr	585F	22623
x"00",	-- Hex Addr	5860	22624
x"00",	-- Hex Addr	5861	22625
x"00",	-- Hex Addr	5862	22626
x"00",	-- Hex Addr	5863	22627
x"00",	-- Hex Addr	5864	22628
x"00",	-- Hex Addr	5865	22629
x"00",	-- Hex Addr	5866	22630
x"00",	-- Hex Addr	5867	22631
x"00",	-- Hex Addr	5868	22632
x"00",	-- Hex Addr	5869	22633
x"00",	-- Hex Addr	586A	22634
x"00",	-- Hex Addr	586B	22635
x"00",	-- Hex Addr	586C	22636
x"00",	-- Hex Addr	586D	22637
x"00",	-- Hex Addr	586E	22638
x"00",	-- Hex Addr	586F	22639
x"00",	-- Hex Addr	5870	22640
x"00",	-- Hex Addr	5871	22641
x"00",	-- Hex Addr	5872	22642
x"00",	-- Hex Addr	5873	22643
x"00",	-- Hex Addr	5874	22644
x"00",	-- Hex Addr	5875	22645
x"00",	-- Hex Addr	5876	22646
x"00",	-- Hex Addr	5877	22647
x"00",	-- Hex Addr	5878	22648
x"00",	-- Hex Addr	5879	22649
x"00",	-- Hex Addr	587A	22650
x"00",	-- Hex Addr	587B	22651
x"00",	-- Hex Addr	587C	22652
x"00",	-- Hex Addr	587D	22653
x"00",	-- Hex Addr	587E	22654
x"00",	-- Hex Addr	587F	22655
x"00",	-- Hex Addr	5880	22656
x"00",	-- Hex Addr	5881	22657
x"00",	-- Hex Addr	5882	22658
x"00",	-- Hex Addr	5883	22659
x"00",	-- Hex Addr	5884	22660
x"00",	-- Hex Addr	5885	22661
x"00",	-- Hex Addr	5886	22662
x"00",	-- Hex Addr	5887	22663
x"00",	-- Hex Addr	5888	22664
x"00",	-- Hex Addr	5889	22665
x"00",	-- Hex Addr	588A	22666
x"00",	-- Hex Addr	588B	22667
x"00",	-- Hex Addr	588C	22668
x"00",	-- Hex Addr	588D	22669
x"00",	-- Hex Addr	588E	22670
x"00",	-- Hex Addr	588F	22671
x"00",	-- Hex Addr	5890	22672
x"00",	-- Hex Addr	5891	22673
x"00",	-- Hex Addr	5892	22674
x"00",	-- Hex Addr	5893	22675
x"00",	-- Hex Addr	5894	22676
x"00",	-- Hex Addr	5895	22677
x"00",	-- Hex Addr	5896	22678
x"00",	-- Hex Addr	5897	22679
x"00",	-- Hex Addr	5898	22680
x"00",	-- Hex Addr	5899	22681
x"00",	-- Hex Addr	589A	22682
x"00",	-- Hex Addr	589B	22683
x"00",	-- Hex Addr	589C	22684
x"00",	-- Hex Addr	589D	22685
x"00",	-- Hex Addr	589E	22686
x"00",	-- Hex Addr	589F	22687
x"00",	-- Hex Addr	58A0	22688
x"00",	-- Hex Addr	58A1	22689
x"00",	-- Hex Addr	58A2	22690
x"00",	-- Hex Addr	58A3	22691
x"00",	-- Hex Addr	58A4	22692
x"00",	-- Hex Addr	58A5	22693
x"00",	-- Hex Addr	58A6	22694
x"00",	-- Hex Addr	58A7	22695
x"00",	-- Hex Addr	58A8	22696
x"00",	-- Hex Addr	58A9	22697
x"00",	-- Hex Addr	58AA	22698
x"00",	-- Hex Addr	58AB	22699
x"00",	-- Hex Addr	58AC	22700
x"00",	-- Hex Addr	58AD	22701
x"00",	-- Hex Addr	58AE	22702
x"00",	-- Hex Addr	58AF	22703
x"00",	-- Hex Addr	58B0	22704
x"00",	-- Hex Addr	58B1	22705
x"00",	-- Hex Addr	58B2	22706
x"00",	-- Hex Addr	58B3	22707
x"00",	-- Hex Addr	58B4	22708
x"00",	-- Hex Addr	58B5	22709
x"00",	-- Hex Addr	58B6	22710
x"00",	-- Hex Addr	58B7	22711
x"00",	-- Hex Addr	58B8	22712
x"00",	-- Hex Addr	58B9	22713
x"00",	-- Hex Addr	58BA	22714
x"00",	-- Hex Addr	58BB	22715
x"00",	-- Hex Addr	58BC	22716
x"00",	-- Hex Addr	58BD	22717
x"00",	-- Hex Addr	58BE	22718
x"00",	-- Hex Addr	58BF	22719
x"00",	-- Hex Addr	58C0	22720
x"00",	-- Hex Addr	58C1	22721
x"00",	-- Hex Addr	58C2	22722
x"00",	-- Hex Addr	58C3	22723
x"00",	-- Hex Addr	58C4	22724
x"00",	-- Hex Addr	58C5	22725
x"00",	-- Hex Addr	58C6	22726
x"00",	-- Hex Addr	58C7	22727
x"00",	-- Hex Addr	58C8	22728
x"00",	-- Hex Addr	58C9	22729
x"00",	-- Hex Addr	58CA	22730
x"00",	-- Hex Addr	58CB	22731
x"00",	-- Hex Addr	58CC	22732
x"00",	-- Hex Addr	58CD	22733
x"00",	-- Hex Addr	58CE	22734
x"00",	-- Hex Addr	58CF	22735
x"00",	-- Hex Addr	58D0	22736
x"00",	-- Hex Addr	58D1	22737
x"00",	-- Hex Addr	58D2	22738
x"00",	-- Hex Addr	58D3	22739
x"00",	-- Hex Addr	58D4	22740
x"00",	-- Hex Addr	58D5	22741
x"00",	-- Hex Addr	58D6	22742
x"00",	-- Hex Addr	58D7	22743
x"00",	-- Hex Addr	58D8	22744
x"00",	-- Hex Addr	58D9	22745
x"00",	-- Hex Addr	58DA	22746
x"00",	-- Hex Addr	58DB	22747
x"00",	-- Hex Addr	58DC	22748
x"00",	-- Hex Addr	58DD	22749
x"00",	-- Hex Addr	58DE	22750
x"00",	-- Hex Addr	58DF	22751
x"00",	-- Hex Addr	58E0	22752
x"00",	-- Hex Addr	58E1	22753
x"00",	-- Hex Addr	58E2	22754
x"00",	-- Hex Addr	58E3	22755
x"00",	-- Hex Addr	58E4	22756
x"00",	-- Hex Addr	58E5	22757
x"00",	-- Hex Addr	58E6	22758
x"00",	-- Hex Addr	58E7	22759
x"00",	-- Hex Addr	58E8	22760
x"00",	-- Hex Addr	58E9	22761
x"00",	-- Hex Addr	58EA	22762
x"00",	-- Hex Addr	58EB	22763
x"00",	-- Hex Addr	58EC	22764
x"00",	-- Hex Addr	58ED	22765
x"00",	-- Hex Addr	58EE	22766
x"00",	-- Hex Addr	58EF	22767
x"00",	-- Hex Addr	58F0	22768
x"00",	-- Hex Addr	58F1	22769
x"00",	-- Hex Addr	58F2	22770
x"00",	-- Hex Addr	58F3	22771
x"00",	-- Hex Addr	58F4	22772
x"00",	-- Hex Addr	58F5	22773
x"00",	-- Hex Addr	58F6	22774
x"00",	-- Hex Addr	58F7	22775
x"00",	-- Hex Addr	58F8	22776
x"00",	-- Hex Addr	58F9	22777
x"00",	-- Hex Addr	58FA	22778
x"00",	-- Hex Addr	58FB	22779
x"00",	-- Hex Addr	58FC	22780
x"00",	-- Hex Addr	58FD	22781
x"00",	-- Hex Addr	58FE	22782
x"00",	-- Hex Addr	58FF	22783
x"00",	-- Hex Addr	5900	22784
x"00",	-- Hex Addr	5901	22785
x"00",	-- Hex Addr	5902	22786
x"00",	-- Hex Addr	5903	22787
x"00",	-- Hex Addr	5904	22788
x"00",	-- Hex Addr	5905	22789
x"00",	-- Hex Addr	5906	22790
x"00",	-- Hex Addr	5907	22791
x"00",	-- Hex Addr	5908	22792
x"00",	-- Hex Addr	5909	22793
x"00",	-- Hex Addr	590A	22794
x"00",	-- Hex Addr	590B	22795
x"00",	-- Hex Addr	590C	22796
x"00",	-- Hex Addr	590D	22797
x"00",	-- Hex Addr	590E	22798
x"00",	-- Hex Addr	590F	22799
x"00",	-- Hex Addr	5910	22800
x"00",	-- Hex Addr	5911	22801
x"00",	-- Hex Addr	5912	22802
x"00",	-- Hex Addr	5913	22803
x"00",	-- Hex Addr	5914	22804
x"00",	-- Hex Addr	5915	22805
x"00",	-- Hex Addr	5916	22806
x"00",	-- Hex Addr	5917	22807
x"00",	-- Hex Addr	5918	22808
x"00",	-- Hex Addr	5919	22809
x"00",	-- Hex Addr	591A	22810
x"00",	-- Hex Addr	591B	22811
x"00",	-- Hex Addr	591C	22812
x"00",	-- Hex Addr	591D	22813
x"00",	-- Hex Addr	591E	22814
x"00",	-- Hex Addr	591F	22815
x"00",	-- Hex Addr	5920	22816
x"00",	-- Hex Addr	5921	22817
x"00",	-- Hex Addr	5922	22818
x"00",	-- Hex Addr	5923	22819
x"00",	-- Hex Addr	5924	22820
x"00",	-- Hex Addr	5925	22821
x"00",	-- Hex Addr	5926	22822
x"00",	-- Hex Addr	5927	22823
x"00",	-- Hex Addr	5928	22824
x"00",	-- Hex Addr	5929	22825
x"00",	-- Hex Addr	592A	22826
x"00",	-- Hex Addr	592B	22827
x"00",	-- Hex Addr	592C	22828
x"00",	-- Hex Addr	592D	22829
x"00",	-- Hex Addr	592E	22830
x"00",	-- Hex Addr	592F	22831
x"00",	-- Hex Addr	5930	22832
x"00",	-- Hex Addr	5931	22833
x"00",	-- Hex Addr	5932	22834
x"00",	-- Hex Addr	5933	22835
x"00",	-- Hex Addr	5934	22836
x"00",	-- Hex Addr	5935	22837
x"00",	-- Hex Addr	5936	22838
x"00",	-- Hex Addr	5937	22839
x"00",	-- Hex Addr	5938	22840
x"00",	-- Hex Addr	5939	22841
x"00",	-- Hex Addr	593A	22842
x"00",	-- Hex Addr	593B	22843
x"00",	-- Hex Addr	593C	22844
x"00",	-- Hex Addr	593D	22845
x"00",	-- Hex Addr	593E	22846
x"00",	-- Hex Addr	593F	22847
x"00",	-- Hex Addr	5940	22848
x"00",	-- Hex Addr	5941	22849
x"00",	-- Hex Addr	5942	22850
x"00",	-- Hex Addr	5943	22851
x"00",	-- Hex Addr	5944	22852
x"00",	-- Hex Addr	5945	22853
x"00",	-- Hex Addr	5946	22854
x"00",	-- Hex Addr	5947	22855
x"00",	-- Hex Addr	5948	22856
x"00",	-- Hex Addr	5949	22857
x"00",	-- Hex Addr	594A	22858
x"00",	-- Hex Addr	594B	22859
x"00",	-- Hex Addr	594C	22860
x"00",	-- Hex Addr	594D	22861
x"00",	-- Hex Addr	594E	22862
x"00",	-- Hex Addr	594F	22863
x"00",	-- Hex Addr	5950	22864
x"00",	-- Hex Addr	5951	22865
x"00",	-- Hex Addr	5952	22866
x"00",	-- Hex Addr	5953	22867
x"00",	-- Hex Addr	5954	22868
x"00",	-- Hex Addr	5955	22869
x"00",	-- Hex Addr	5956	22870
x"00",	-- Hex Addr	5957	22871
x"00",	-- Hex Addr	5958	22872
x"00",	-- Hex Addr	5959	22873
x"00",	-- Hex Addr	595A	22874
x"00",	-- Hex Addr	595B	22875
x"00",	-- Hex Addr	595C	22876
x"00",	-- Hex Addr	595D	22877
x"00",	-- Hex Addr	595E	22878
x"00",	-- Hex Addr	595F	22879
x"00",	-- Hex Addr	5960	22880
x"00",	-- Hex Addr	5961	22881
x"00",	-- Hex Addr	5962	22882
x"00",	-- Hex Addr	5963	22883
x"00",	-- Hex Addr	5964	22884
x"00",	-- Hex Addr	5965	22885
x"00",	-- Hex Addr	5966	22886
x"00",	-- Hex Addr	5967	22887
x"00",	-- Hex Addr	5968	22888
x"00",	-- Hex Addr	5969	22889
x"00",	-- Hex Addr	596A	22890
x"00",	-- Hex Addr	596B	22891
x"00",	-- Hex Addr	596C	22892
x"00",	-- Hex Addr	596D	22893
x"00",	-- Hex Addr	596E	22894
x"00",	-- Hex Addr	596F	22895
x"00",	-- Hex Addr	5970	22896
x"00",	-- Hex Addr	5971	22897
x"00",	-- Hex Addr	5972	22898
x"00",	-- Hex Addr	5973	22899
x"00",	-- Hex Addr	5974	22900
x"00",	-- Hex Addr	5975	22901
x"00",	-- Hex Addr	5976	22902
x"00",	-- Hex Addr	5977	22903
x"00",	-- Hex Addr	5978	22904
x"00",	-- Hex Addr	5979	22905
x"00",	-- Hex Addr	597A	22906
x"00",	-- Hex Addr	597B	22907
x"00",	-- Hex Addr	597C	22908
x"00",	-- Hex Addr	597D	22909
x"00",	-- Hex Addr	597E	22910
x"00",	-- Hex Addr	597F	22911
x"00",	-- Hex Addr	5980	22912
x"00",	-- Hex Addr	5981	22913
x"00",	-- Hex Addr	5982	22914
x"00",	-- Hex Addr	5983	22915
x"00",	-- Hex Addr	5984	22916
x"00",	-- Hex Addr	5985	22917
x"00",	-- Hex Addr	5986	22918
x"00",	-- Hex Addr	5987	22919
x"00",	-- Hex Addr	5988	22920
x"00",	-- Hex Addr	5989	22921
x"00",	-- Hex Addr	598A	22922
x"00",	-- Hex Addr	598B	22923
x"00",	-- Hex Addr	598C	22924
x"00",	-- Hex Addr	598D	22925
x"00",	-- Hex Addr	598E	22926
x"00",	-- Hex Addr	598F	22927
x"00",	-- Hex Addr	5990	22928
x"00",	-- Hex Addr	5991	22929
x"00",	-- Hex Addr	5992	22930
x"00",	-- Hex Addr	5993	22931
x"00",	-- Hex Addr	5994	22932
x"00",	-- Hex Addr	5995	22933
x"00",	-- Hex Addr	5996	22934
x"00",	-- Hex Addr	5997	22935
x"00",	-- Hex Addr	5998	22936
x"00",	-- Hex Addr	5999	22937
x"00",	-- Hex Addr	599A	22938
x"00",	-- Hex Addr	599B	22939
x"00",	-- Hex Addr	599C	22940
x"00",	-- Hex Addr	599D	22941
x"00",	-- Hex Addr	599E	22942
x"00",	-- Hex Addr	599F	22943
x"00",	-- Hex Addr	59A0	22944
x"00",	-- Hex Addr	59A1	22945
x"00",	-- Hex Addr	59A2	22946
x"00",	-- Hex Addr	59A3	22947
x"00",	-- Hex Addr	59A4	22948
x"00",	-- Hex Addr	59A5	22949
x"00",	-- Hex Addr	59A6	22950
x"00",	-- Hex Addr	59A7	22951
x"00",	-- Hex Addr	59A8	22952
x"00",	-- Hex Addr	59A9	22953
x"00",	-- Hex Addr	59AA	22954
x"00",	-- Hex Addr	59AB	22955
x"00",	-- Hex Addr	59AC	22956
x"00",	-- Hex Addr	59AD	22957
x"00",	-- Hex Addr	59AE	22958
x"00",	-- Hex Addr	59AF	22959
x"00",	-- Hex Addr	59B0	22960
x"00",	-- Hex Addr	59B1	22961
x"00",	-- Hex Addr	59B2	22962
x"00",	-- Hex Addr	59B3	22963
x"00",	-- Hex Addr	59B4	22964
x"00",	-- Hex Addr	59B5	22965
x"00",	-- Hex Addr	59B6	22966
x"00",	-- Hex Addr	59B7	22967
x"00",	-- Hex Addr	59B8	22968
x"00",	-- Hex Addr	59B9	22969
x"00",	-- Hex Addr	59BA	22970
x"00",	-- Hex Addr	59BB	22971
x"00",	-- Hex Addr	59BC	22972
x"00",	-- Hex Addr	59BD	22973
x"00",	-- Hex Addr	59BE	22974
x"00",	-- Hex Addr	59BF	22975
x"00",	-- Hex Addr	59C0	22976
x"00",	-- Hex Addr	59C1	22977
x"00",	-- Hex Addr	59C2	22978
x"00",	-- Hex Addr	59C3	22979
x"00",	-- Hex Addr	59C4	22980
x"00",	-- Hex Addr	59C5	22981
x"00",	-- Hex Addr	59C6	22982
x"00",	-- Hex Addr	59C7	22983
x"00",	-- Hex Addr	59C8	22984
x"00",	-- Hex Addr	59C9	22985
x"00",	-- Hex Addr	59CA	22986
x"00",	-- Hex Addr	59CB	22987
x"00",	-- Hex Addr	59CC	22988
x"00",	-- Hex Addr	59CD	22989
x"00",	-- Hex Addr	59CE	22990
x"00",	-- Hex Addr	59CF	22991
x"00",	-- Hex Addr	59D0	22992
x"00",	-- Hex Addr	59D1	22993
x"00",	-- Hex Addr	59D2	22994
x"00",	-- Hex Addr	59D3	22995
x"00",	-- Hex Addr	59D4	22996
x"00",	-- Hex Addr	59D5	22997
x"00",	-- Hex Addr	59D6	22998
x"00",	-- Hex Addr	59D7	22999
x"00",	-- Hex Addr	59D8	23000
x"00",	-- Hex Addr	59D9	23001
x"00",	-- Hex Addr	59DA	23002
x"00",	-- Hex Addr	59DB	23003
x"00",	-- Hex Addr	59DC	23004
x"00",	-- Hex Addr	59DD	23005
x"00",	-- Hex Addr	59DE	23006
x"00",	-- Hex Addr	59DF	23007
x"00",	-- Hex Addr	59E0	23008
x"00",	-- Hex Addr	59E1	23009
x"00",	-- Hex Addr	59E2	23010
x"00",	-- Hex Addr	59E3	23011
x"00",	-- Hex Addr	59E4	23012
x"00",	-- Hex Addr	59E5	23013
x"00",	-- Hex Addr	59E6	23014
x"00",	-- Hex Addr	59E7	23015
x"00",	-- Hex Addr	59E8	23016
x"00",	-- Hex Addr	59E9	23017
x"00",	-- Hex Addr	59EA	23018
x"00",	-- Hex Addr	59EB	23019
x"00",	-- Hex Addr	59EC	23020
x"00",	-- Hex Addr	59ED	23021
x"00",	-- Hex Addr	59EE	23022
x"00",	-- Hex Addr	59EF	23023
x"00",	-- Hex Addr	59F0	23024
x"00",	-- Hex Addr	59F1	23025
x"00",	-- Hex Addr	59F2	23026
x"00",	-- Hex Addr	59F3	23027
x"00",	-- Hex Addr	59F4	23028
x"00",	-- Hex Addr	59F5	23029
x"00",	-- Hex Addr	59F6	23030
x"00",	-- Hex Addr	59F7	23031
x"00",	-- Hex Addr	59F8	23032
x"00",	-- Hex Addr	59F9	23033
x"00",	-- Hex Addr	59FA	23034
x"00",	-- Hex Addr	59FB	23035
x"00",	-- Hex Addr	59FC	23036
x"00",	-- Hex Addr	59FD	23037
x"00",	-- Hex Addr	59FE	23038
x"00",	-- Hex Addr	59FF	23039
x"00",	-- Hex Addr	5A00	23040
x"00",	-- Hex Addr	5A01	23041
x"00",	-- Hex Addr	5A02	23042
x"00",	-- Hex Addr	5A03	23043
x"00",	-- Hex Addr	5A04	23044
x"00",	-- Hex Addr	5A05	23045
x"00",	-- Hex Addr	5A06	23046
x"00",	-- Hex Addr	5A07	23047
x"00",	-- Hex Addr	5A08	23048
x"00",	-- Hex Addr	5A09	23049
x"00",	-- Hex Addr	5A0A	23050
x"00",	-- Hex Addr	5A0B	23051
x"00",	-- Hex Addr	5A0C	23052
x"00",	-- Hex Addr	5A0D	23053
x"00",	-- Hex Addr	5A0E	23054
x"00",	-- Hex Addr	5A0F	23055
x"00",	-- Hex Addr	5A10	23056
x"00",	-- Hex Addr	5A11	23057
x"00",	-- Hex Addr	5A12	23058
x"00",	-- Hex Addr	5A13	23059
x"00",	-- Hex Addr	5A14	23060
x"00",	-- Hex Addr	5A15	23061
x"00",	-- Hex Addr	5A16	23062
x"00",	-- Hex Addr	5A17	23063
x"00",	-- Hex Addr	5A18	23064
x"00",	-- Hex Addr	5A19	23065
x"00",	-- Hex Addr	5A1A	23066
x"00",	-- Hex Addr	5A1B	23067
x"00",	-- Hex Addr	5A1C	23068
x"00",	-- Hex Addr	5A1D	23069
x"00",	-- Hex Addr	5A1E	23070
x"00",	-- Hex Addr	5A1F	23071
x"00",	-- Hex Addr	5A20	23072
x"00",	-- Hex Addr	5A21	23073
x"00",	-- Hex Addr	5A22	23074
x"00",	-- Hex Addr	5A23	23075
x"00",	-- Hex Addr	5A24	23076
x"00",	-- Hex Addr	5A25	23077
x"00",	-- Hex Addr	5A26	23078
x"00",	-- Hex Addr	5A27	23079
x"00",	-- Hex Addr	5A28	23080
x"00",	-- Hex Addr	5A29	23081
x"00",	-- Hex Addr	5A2A	23082
x"00",	-- Hex Addr	5A2B	23083
x"00",	-- Hex Addr	5A2C	23084
x"00",	-- Hex Addr	5A2D	23085
x"00",	-- Hex Addr	5A2E	23086
x"00",	-- Hex Addr	5A2F	23087
x"00",	-- Hex Addr	5A30	23088
x"00",	-- Hex Addr	5A31	23089
x"00",	-- Hex Addr	5A32	23090
x"00",	-- Hex Addr	5A33	23091
x"00",	-- Hex Addr	5A34	23092
x"00",	-- Hex Addr	5A35	23093
x"00",	-- Hex Addr	5A36	23094
x"00",	-- Hex Addr	5A37	23095
x"00",	-- Hex Addr	5A38	23096
x"00",	-- Hex Addr	5A39	23097
x"00",	-- Hex Addr	5A3A	23098
x"00",	-- Hex Addr	5A3B	23099
x"00",	-- Hex Addr	5A3C	23100
x"00",	-- Hex Addr	5A3D	23101
x"00",	-- Hex Addr	5A3E	23102
x"00",	-- Hex Addr	5A3F	23103
x"00",	-- Hex Addr	5A40	23104
x"00",	-- Hex Addr	5A41	23105
x"00",	-- Hex Addr	5A42	23106
x"00",	-- Hex Addr	5A43	23107
x"00",	-- Hex Addr	5A44	23108
x"00",	-- Hex Addr	5A45	23109
x"00",	-- Hex Addr	5A46	23110
x"00",	-- Hex Addr	5A47	23111
x"00",	-- Hex Addr	5A48	23112
x"00",	-- Hex Addr	5A49	23113
x"00",	-- Hex Addr	5A4A	23114
x"00",	-- Hex Addr	5A4B	23115
x"00",	-- Hex Addr	5A4C	23116
x"00",	-- Hex Addr	5A4D	23117
x"00",	-- Hex Addr	5A4E	23118
x"00",	-- Hex Addr	5A4F	23119
x"00",	-- Hex Addr	5A50	23120
x"00",	-- Hex Addr	5A51	23121
x"00",	-- Hex Addr	5A52	23122
x"00",	-- Hex Addr	5A53	23123
x"00",	-- Hex Addr	5A54	23124
x"00",	-- Hex Addr	5A55	23125
x"00",	-- Hex Addr	5A56	23126
x"00",	-- Hex Addr	5A57	23127
x"00",	-- Hex Addr	5A58	23128
x"00",	-- Hex Addr	5A59	23129
x"00",	-- Hex Addr	5A5A	23130
x"00",	-- Hex Addr	5A5B	23131
x"00",	-- Hex Addr	5A5C	23132
x"00",	-- Hex Addr	5A5D	23133
x"00",	-- Hex Addr	5A5E	23134
x"00",	-- Hex Addr	5A5F	23135
x"00",	-- Hex Addr	5A60	23136
x"00",	-- Hex Addr	5A61	23137
x"00",	-- Hex Addr	5A62	23138
x"00",	-- Hex Addr	5A63	23139
x"00",	-- Hex Addr	5A64	23140
x"00",	-- Hex Addr	5A65	23141
x"00",	-- Hex Addr	5A66	23142
x"00",	-- Hex Addr	5A67	23143
x"00",	-- Hex Addr	5A68	23144
x"00",	-- Hex Addr	5A69	23145
x"00",	-- Hex Addr	5A6A	23146
x"00",	-- Hex Addr	5A6B	23147
x"00",	-- Hex Addr	5A6C	23148
x"00",	-- Hex Addr	5A6D	23149
x"00",	-- Hex Addr	5A6E	23150
x"00",	-- Hex Addr	5A6F	23151
x"00",	-- Hex Addr	5A70	23152
x"00",	-- Hex Addr	5A71	23153
x"00",	-- Hex Addr	5A72	23154
x"00",	-- Hex Addr	5A73	23155
x"00",	-- Hex Addr	5A74	23156
x"00",	-- Hex Addr	5A75	23157
x"00",	-- Hex Addr	5A76	23158
x"00",	-- Hex Addr	5A77	23159
x"00",	-- Hex Addr	5A78	23160
x"00",	-- Hex Addr	5A79	23161
x"00",	-- Hex Addr	5A7A	23162
x"00",	-- Hex Addr	5A7B	23163
x"00",	-- Hex Addr	5A7C	23164
x"00",	-- Hex Addr	5A7D	23165
x"00",	-- Hex Addr	5A7E	23166
x"00",	-- Hex Addr	5A7F	23167
x"00",	-- Hex Addr	5A80	23168
x"00",	-- Hex Addr	5A81	23169
x"00",	-- Hex Addr	5A82	23170
x"00",	-- Hex Addr	5A83	23171
x"00",	-- Hex Addr	5A84	23172
x"00",	-- Hex Addr	5A85	23173
x"00",	-- Hex Addr	5A86	23174
x"00",	-- Hex Addr	5A87	23175
x"00",	-- Hex Addr	5A88	23176
x"00",	-- Hex Addr	5A89	23177
x"00",	-- Hex Addr	5A8A	23178
x"00",	-- Hex Addr	5A8B	23179
x"00",	-- Hex Addr	5A8C	23180
x"00",	-- Hex Addr	5A8D	23181
x"00",	-- Hex Addr	5A8E	23182
x"00",	-- Hex Addr	5A8F	23183
x"00",	-- Hex Addr	5A90	23184
x"00",	-- Hex Addr	5A91	23185
x"00",	-- Hex Addr	5A92	23186
x"00",	-- Hex Addr	5A93	23187
x"00",	-- Hex Addr	5A94	23188
x"00",	-- Hex Addr	5A95	23189
x"00",	-- Hex Addr	5A96	23190
x"00",	-- Hex Addr	5A97	23191
x"00",	-- Hex Addr	5A98	23192
x"00",	-- Hex Addr	5A99	23193
x"00",	-- Hex Addr	5A9A	23194
x"00",	-- Hex Addr	5A9B	23195
x"00",	-- Hex Addr	5A9C	23196
x"00",	-- Hex Addr	5A9D	23197
x"00",	-- Hex Addr	5A9E	23198
x"00",	-- Hex Addr	5A9F	23199
x"00",	-- Hex Addr	5AA0	23200
x"00",	-- Hex Addr	5AA1	23201
x"00",	-- Hex Addr	5AA2	23202
x"00",	-- Hex Addr	5AA3	23203
x"00",	-- Hex Addr	5AA4	23204
x"00",	-- Hex Addr	5AA5	23205
x"00",	-- Hex Addr	5AA6	23206
x"00",	-- Hex Addr	5AA7	23207
x"00",	-- Hex Addr	5AA8	23208
x"00",	-- Hex Addr	5AA9	23209
x"00",	-- Hex Addr	5AAA	23210
x"00",	-- Hex Addr	5AAB	23211
x"00",	-- Hex Addr	5AAC	23212
x"00",	-- Hex Addr	5AAD	23213
x"00",	-- Hex Addr	5AAE	23214
x"00",	-- Hex Addr	5AAF	23215
x"00",	-- Hex Addr	5AB0	23216
x"00",	-- Hex Addr	5AB1	23217
x"00",	-- Hex Addr	5AB2	23218
x"00",	-- Hex Addr	5AB3	23219
x"00",	-- Hex Addr	5AB4	23220
x"00",	-- Hex Addr	5AB5	23221
x"00",	-- Hex Addr	5AB6	23222
x"00",	-- Hex Addr	5AB7	23223
x"00",	-- Hex Addr	5AB8	23224
x"00",	-- Hex Addr	5AB9	23225
x"00",	-- Hex Addr	5ABA	23226
x"00",	-- Hex Addr	5ABB	23227
x"00",	-- Hex Addr	5ABC	23228
x"00",	-- Hex Addr	5ABD	23229
x"00",	-- Hex Addr	5ABE	23230
x"00",	-- Hex Addr	5ABF	23231
x"00",	-- Hex Addr	5AC0	23232
x"00",	-- Hex Addr	5AC1	23233
x"00",	-- Hex Addr	5AC2	23234
x"00",	-- Hex Addr	5AC3	23235
x"00",	-- Hex Addr	5AC4	23236
x"00",	-- Hex Addr	5AC5	23237
x"00",	-- Hex Addr	5AC6	23238
x"00",	-- Hex Addr	5AC7	23239
x"00",	-- Hex Addr	5AC8	23240
x"00",	-- Hex Addr	5AC9	23241
x"00",	-- Hex Addr	5ACA	23242
x"00",	-- Hex Addr	5ACB	23243
x"00",	-- Hex Addr	5ACC	23244
x"00",	-- Hex Addr	5ACD	23245
x"00",	-- Hex Addr	5ACE	23246
x"00",	-- Hex Addr	5ACF	23247
x"00",	-- Hex Addr	5AD0	23248
x"00",	-- Hex Addr	5AD1	23249
x"00",	-- Hex Addr	5AD2	23250
x"00",	-- Hex Addr	5AD3	23251
x"00",	-- Hex Addr	5AD4	23252
x"00",	-- Hex Addr	5AD5	23253
x"00",	-- Hex Addr	5AD6	23254
x"00",	-- Hex Addr	5AD7	23255
x"00",	-- Hex Addr	5AD8	23256
x"00",	-- Hex Addr	5AD9	23257
x"00",	-- Hex Addr	5ADA	23258
x"00",	-- Hex Addr	5ADB	23259
x"00",	-- Hex Addr	5ADC	23260
x"00",	-- Hex Addr	5ADD	23261
x"00",	-- Hex Addr	5ADE	23262
x"00",	-- Hex Addr	5ADF	23263
x"00",	-- Hex Addr	5AE0	23264
x"00",	-- Hex Addr	5AE1	23265
x"00",	-- Hex Addr	5AE2	23266
x"00",	-- Hex Addr	5AE3	23267
x"00",	-- Hex Addr	5AE4	23268
x"00",	-- Hex Addr	5AE5	23269
x"00",	-- Hex Addr	5AE6	23270
x"00",	-- Hex Addr	5AE7	23271
x"00",	-- Hex Addr	5AE8	23272
x"00",	-- Hex Addr	5AE9	23273
x"00",	-- Hex Addr	5AEA	23274
x"00",	-- Hex Addr	5AEB	23275
x"00",	-- Hex Addr	5AEC	23276
x"00",	-- Hex Addr	5AED	23277
x"00",	-- Hex Addr	5AEE	23278
x"00",	-- Hex Addr	5AEF	23279
x"00",	-- Hex Addr	5AF0	23280
x"00",	-- Hex Addr	5AF1	23281
x"00",	-- Hex Addr	5AF2	23282
x"00",	-- Hex Addr	5AF3	23283
x"00",	-- Hex Addr	5AF4	23284
x"00",	-- Hex Addr	5AF5	23285
x"00",	-- Hex Addr	5AF6	23286
x"00",	-- Hex Addr	5AF7	23287
x"00",	-- Hex Addr	5AF8	23288
x"00",	-- Hex Addr	5AF9	23289
x"00",	-- Hex Addr	5AFA	23290
x"00",	-- Hex Addr	5AFB	23291
x"00",	-- Hex Addr	5AFC	23292
x"00",	-- Hex Addr	5AFD	23293
x"00",	-- Hex Addr	5AFE	23294
x"00",	-- Hex Addr	5AFF	23295
x"00",	-- Hex Addr	5B00	23296
x"00",	-- Hex Addr	5B01	23297
x"00",	-- Hex Addr	5B02	23298
x"00",	-- Hex Addr	5B03	23299
x"00",	-- Hex Addr	5B04	23300
x"00",	-- Hex Addr	5B05	23301
x"00",	-- Hex Addr	5B06	23302
x"00",	-- Hex Addr	5B07	23303
x"00",	-- Hex Addr	5B08	23304
x"00",	-- Hex Addr	5B09	23305
x"00",	-- Hex Addr	5B0A	23306
x"00",	-- Hex Addr	5B0B	23307
x"00",	-- Hex Addr	5B0C	23308
x"00",	-- Hex Addr	5B0D	23309
x"00",	-- Hex Addr	5B0E	23310
x"00",	-- Hex Addr	5B0F	23311
x"00",	-- Hex Addr	5B10	23312
x"00",	-- Hex Addr	5B11	23313
x"00",	-- Hex Addr	5B12	23314
x"00",	-- Hex Addr	5B13	23315
x"00",	-- Hex Addr	5B14	23316
x"00",	-- Hex Addr	5B15	23317
x"00",	-- Hex Addr	5B16	23318
x"00",	-- Hex Addr	5B17	23319
x"00",	-- Hex Addr	5B18	23320
x"00",	-- Hex Addr	5B19	23321
x"00",	-- Hex Addr	5B1A	23322
x"00",	-- Hex Addr	5B1B	23323
x"00",	-- Hex Addr	5B1C	23324
x"00",	-- Hex Addr	5B1D	23325
x"00",	-- Hex Addr	5B1E	23326
x"00",	-- Hex Addr	5B1F	23327
x"00",	-- Hex Addr	5B20	23328
x"00",	-- Hex Addr	5B21	23329
x"00",	-- Hex Addr	5B22	23330
x"00",	-- Hex Addr	5B23	23331
x"00",	-- Hex Addr	5B24	23332
x"00",	-- Hex Addr	5B25	23333
x"00",	-- Hex Addr	5B26	23334
x"00",	-- Hex Addr	5B27	23335
x"00",	-- Hex Addr	5B28	23336
x"00",	-- Hex Addr	5B29	23337
x"00",	-- Hex Addr	5B2A	23338
x"00",	-- Hex Addr	5B2B	23339
x"00",	-- Hex Addr	5B2C	23340
x"00",	-- Hex Addr	5B2D	23341
x"00",	-- Hex Addr	5B2E	23342
x"00",	-- Hex Addr	5B2F	23343
x"00",	-- Hex Addr	5B30	23344
x"00",	-- Hex Addr	5B31	23345
x"00",	-- Hex Addr	5B32	23346
x"00",	-- Hex Addr	5B33	23347
x"00",	-- Hex Addr	5B34	23348
x"00",	-- Hex Addr	5B35	23349
x"00",	-- Hex Addr	5B36	23350
x"00",	-- Hex Addr	5B37	23351
x"00",	-- Hex Addr	5B38	23352
x"00",	-- Hex Addr	5B39	23353
x"00",	-- Hex Addr	5B3A	23354
x"00",	-- Hex Addr	5B3B	23355
x"00",	-- Hex Addr	5B3C	23356
x"00",	-- Hex Addr	5B3D	23357
x"00",	-- Hex Addr	5B3E	23358
x"00",	-- Hex Addr	5B3F	23359
x"00",	-- Hex Addr	5B40	23360
x"00",	-- Hex Addr	5B41	23361
x"00",	-- Hex Addr	5B42	23362
x"00",	-- Hex Addr	5B43	23363
x"00",	-- Hex Addr	5B44	23364
x"00",	-- Hex Addr	5B45	23365
x"00",	-- Hex Addr	5B46	23366
x"00",	-- Hex Addr	5B47	23367
x"00",	-- Hex Addr	5B48	23368
x"00",	-- Hex Addr	5B49	23369
x"00",	-- Hex Addr	5B4A	23370
x"00",	-- Hex Addr	5B4B	23371
x"00",	-- Hex Addr	5B4C	23372
x"00",	-- Hex Addr	5B4D	23373
x"00",	-- Hex Addr	5B4E	23374
x"00",	-- Hex Addr	5B4F	23375
x"00",	-- Hex Addr	5B50	23376
x"00",	-- Hex Addr	5B51	23377
x"00",	-- Hex Addr	5B52	23378
x"00",	-- Hex Addr	5B53	23379
x"00",	-- Hex Addr	5B54	23380
x"00",	-- Hex Addr	5B55	23381
x"00",	-- Hex Addr	5B56	23382
x"00",	-- Hex Addr	5B57	23383
x"00",	-- Hex Addr	5B58	23384
x"00",	-- Hex Addr	5B59	23385
x"00",	-- Hex Addr	5B5A	23386
x"00",	-- Hex Addr	5B5B	23387
x"00",	-- Hex Addr	5B5C	23388
x"00",	-- Hex Addr	5B5D	23389
x"00",	-- Hex Addr	5B5E	23390
x"00",	-- Hex Addr	5B5F	23391
x"00",	-- Hex Addr	5B60	23392
x"00",	-- Hex Addr	5B61	23393
x"00",	-- Hex Addr	5B62	23394
x"00",	-- Hex Addr	5B63	23395
x"00",	-- Hex Addr	5B64	23396
x"00",	-- Hex Addr	5B65	23397
x"00",	-- Hex Addr	5B66	23398
x"00",	-- Hex Addr	5B67	23399
x"00",	-- Hex Addr	5B68	23400
x"00",	-- Hex Addr	5B69	23401
x"00",	-- Hex Addr	5B6A	23402
x"00",	-- Hex Addr	5B6B	23403
x"00",	-- Hex Addr	5B6C	23404
x"00",	-- Hex Addr	5B6D	23405
x"00",	-- Hex Addr	5B6E	23406
x"00",	-- Hex Addr	5B6F	23407
x"00",	-- Hex Addr	5B70	23408
x"00",	-- Hex Addr	5B71	23409
x"00",	-- Hex Addr	5B72	23410
x"00",	-- Hex Addr	5B73	23411
x"00",	-- Hex Addr	5B74	23412
x"00",	-- Hex Addr	5B75	23413
x"00",	-- Hex Addr	5B76	23414
x"00",	-- Hex Addr	5B77	23415
x"00",	-- Hex Addr	5B78	23416
x"00",	-- Hex Addr	5B79	23417
x"00",	-- Hex Addr	5B7A	23418
x"00",	-- Hex Addr	5B7B	23419
x"00",	-- Hex Addr	5B7C	23420
x"00",	-- Hex Addr	5B7D	23421
x"00",	-- Hex Addr	5B7E	23422
x"00",	-- Hex Addr	5B7F	23423
x"00",	-- Hex Addr	5B80	23424
x"00",	-- Hex Addr	5B81	23425
x"00",	-- Hex Addr	5B82	23426
x"00",	-- Hex Addr	5B83	23427
x"00",	-- Hex Addr	5B84	23428
x"00",	-- Hex Addr	5B85	23429
x"00",	-- Hex Addr	5B86	23430
x"00",	-- Hex Addr	5B87	23431
x"00",	-- Hex Addr	5B88	23432
x"00",	-- Hex Addr	5B89	23433
x"00",	-- Hex Addr	5B8A	23434
x"00",	-- Hex Addr	5B8B	23435
x"00",	-- Hex Addr	5B8C	23436
x"00",	-- Hex Addr	5B8D	23437
x"00",	-- Hex Addr	5B8E	23438
x"00",	-- Hex Addr	5B8F	23439
x"00",	-- Hex Addr	5B90	23440
x"00",	-- Hex Addr	5B91	23441
x"00",	-- Hex Addr	5B92	23442
x"00",	-- Hex Addr	5B93	23443
x"00",	-- Hex Addr	5B94	23444
x"00",	-- Hex Addr	5B95	23445
x"00",	-- Hex Addr	5B96	23446
x"00",	-- Hex Addr	5B97	23447
x"00",	-- Hex Addr	5B98	23448
x"00",	-- Hex Addr	5B99	23449
x"00",	-- Hex Addr	5B9A	23450
x"00",	-- Hex Addr	5B9B	23451
x"00",	-- Hex Addr	5B9C	23452
x"00",	-- Hex Addr	5B9D	23453
x"00",	-- Hex Addr	5B9E	23454
x"00",	-- Hex Addr	5B9F	23455
x"00",	-- Hex Addr	5BA0	23456
x"00",	-- Hex Addr	5BA1	23457
x"00",	-- Hex Addr	5BA2	23458
x"00",	-- Hex Addr	5BA3	23459
x"00",	-- Hex Addr	5BA4	23460
x"00",	-- Hex Addr	5BA5	23461
x"00",	-- Hex Addr	5BA6	23462
x"00",	-- Hex Addr	5BA7	23463
x"00",	-- Hex Addr	5BA8	23464
x"00",	-- Hex Addr	5BA9	23465
x"00",	-- Hex Addr	5BAA	23466
x"00",	-- Hex Addr	5BAB	23467
x"00",	-- Hex Addr	5BAC	23468
x"00",	-- Hex Addr	5BAD	23469
x"00",	-- Hex Addr	5BAE	23470
x"00",	-- Hex Addr	5BAF	23471
x"00",	-- Hex Addr	5BB0	23472
x"00",	-- Hex Addr	5BB1	23473
x"00",	-- Hex Addr	5BB2	23474
x"00",	-- Hex Addr	5BB3	23475
x"00",	-- Hex Addr	5BB4	23476
x"00",	-- Hex Addr	5BB5	23477
x"00",	-- Hex Addr	5BB6	23478
x"00",	-- Hex Addr	5BB7	23479
x"00",	-- Hex Addr	5BB8	23480
x"00",	-- Hex Addr	5BB9	23481
x"00",	-- Hex Addr	5BBA	23482
x"00",	-- Hex Addr	5BBB	23483
x"00",	-- Hex Addr	5BBC	23484
x"00",	-- Hex Addr	5BBD	23485
x"00",	-- Hex Addr	5BBE	23486
x"00",	-- Hex Addr	5BBF	23487
x"00",	-- Hex Addr	5BC0	23488
x"00",	-- Hex Addr	5BC1	23489
x"00",	-- Hex Addr	5BC2	23490
x"00",	-- Hex Addr	5BC3	23491
x"00",	-- Hex Addr	5BC4	23492
x"00",	-- Hex Addr	5BC5	23493
x"00",	-- Hex Addr	5BC6	23494
x"00",	-- Hex Addr	5BC7	23495
x"00",	-- Hex Addr	5BC8	23496
x"00",	-- Hex Addr	5BC9	23497
x"00",	-- Hex Addr	5BCA	23498
x"00",	-- Hex Addr	5BCB	23499
x"00",	-- Hex Addr	5BCC	23500
x"00",	-- Hex Addr	5BCD	23501
x"00",	-- Hex Addr	5BCE	23502
x"00",	-- Hex Addr	5BCF	23503
x"00",	-- Hex Addr	5BD0	23504
x"00",	-- Hex Addr	5BD1	23505
x"00",	-- Hex Addr	5BD2	23506
x"00",	-- Hex Addr	5BD3	23507
x"00",	-- Hex Addr	5BD4	23508
x"00",	-- Hex Addr	5BD5	23509
x"00",	-- Hex Addr	5BD6	23510
x"00",	-- Hex Addr	5BD7	23511
x"00",	-- Hex Addr	5BD8	23512
x"00",	-- Hex Addr	5BD9	23513
x"00",	-- Hex Addr	5BDA	23514
x"00",	-- Hex Addr	5BDB	23515
x"00",	-- Hex Addr	5BDC	23516
x"00",	-- Hex Addr	5BDD	23517
x"00",	-- Hex Addr	5BDE	23518
x"00",	-- Hex Addr	5BDF	23519
x"00",	-- Hex Addr	5BE0	23520
x"00",	-- Hex Addr	5BE1	23521
x"00",	-- Hex Addr	5BE2	23522
x"00",	-- Hex Addr	5BE3	23523
x"00",	-- Hex Addr	5BE4	23524
x"00",	-- Hex Addr	5BE5	23525
x"00",	-- Hex Addr	5BE6	23526
x"00",	-- Hex Addr	5BE7	23527
x"00",	-- Hex Addr	5BE8	23528
x"00",	-- Hex Addr	5BE9	23529
x"00",	-- Hex Addr	5BEA	23530
x"00",	-- Hex Addr	5BEB	23531
x"00",	-- Hex Addr	5BEC	23532
x"00",	-- Hex Addr	5BED	23533
x"00",	-- Hex Addr	5BEE	23534
x"00",	-- Hex Addr	5BEF	23535
x"00",	-- Hex Addr	5BF0	23536
x"00",	-- Hex Addr	5BF1	23537
x"00",	-- Hex Addr	5BF2	23538
x"00",	-- Hex Addr	5BF3	23539
x"00",	-- Hex Addr	5BF4	23540
x"00",	-- Hex Addr	5BF5	23541
x"00",	-- Hex Addr	5BF6	23542
x"00",	-- Hex Addr	5BF7	23543
x"00",	-- Hex Addr	5BF8	23544
x"00",	-- Hex Addr	5BF9	23545
x"00",	-- Hex Addr	5BFA	23546
x"00",	-- Hex Addr	5BFB	23547
x"00",	-- Hex Addr	5BFC	23548
x"00",	-- Hex Addr	5BFD	23549
x"00",	-- Hex Addr	5BFE	23550
x"00",	-- Hex Addr	5BFF	23551
x"00",	-- Hex Addr	5C00	23552
x"00",	-- Hex Addr	5C01	23553
x"00",	-- Hex Addr	5C02	23554
x"00",	-- Hex Addr	5C03	23555
x"00",	-- Hex Addr	5C04	23556
x"00",	-- Hex Addr	5C05	23557
x"00",	-- Hex Addr	5C06	23558
x"00",	-- Hex Addr	5C07	23559
x"00",	-- Hex Addr	5C08	23560
x"00",	-- Hex Addr	5C09	23561
x"00",	-- Hex Addr	5C0A	23562
x"00",	-- Hex Addr	5C0B	23563
x"00",	-- Hex Addr	5C0C	23564
x"00",	-- Hex Addr	5C0D	23565
x"00",	-- Hex Addr	5C0E	23566
x"00",	-- Hex Addr	5C0F	23567
x"00",	-- Hex Addr	5C10	23568
x"00",	-- Hex Addr	5C11	23569
x"00",	-- Hex Addr	5C12	23570
x"00",	-- Hex Addr	5C13	23571
x"00",	-- Hex Addr	5C14	23572
x"00",	-- Hex Addr	5C15	23573
x"00",	-- Hex Addr	5C16	23574
x"00",	-- Hex Addr	5C17	23575
x"00",	-- Hex Addr	5C18	23576
x"00",	-- Hex Addr	5C19	23577
x"00",	-- Hex Addr	5C1A	23578
x"00",	-- Hex Addr	5C1B	23579
x"00",	-- Hex Addr	5C1C	23580
x"00",	-- Hex Addr	5C1D	23581
x"00",	-- Hex Addr	5C1E	23582
x"00",	-- Hex Addr	5C1F	23583
x"00",	-- Hex Addr	5C20	23584
x"00",	-- Hex Addr	5C21	23585
x"00",	-- Hex Addr	5C22	23586
x"00",	-- Hex Addr	5C23	23587
x"00",	-- Hex Addr	5C24	23588
x"00",	-- Hex Addr	5C25	23589
x"00",	-- Hex Addr	5C26	23590
x"00",	-- Hex Addr	5C27	23591
x"00",	-- Hex Addr	5C28	23592
x"00",	-- Hex Addr	5C29	23593
x"00",	-- Hex Addr	5C2A	23594
x"00",	-- Hex Addr	5C2B	23595
x"00",	-- Hex Addr	5C2C	23596
x"00",	-- Hex Addr	5C2D	23597
x"00",	-- Hex Addr	5C2E	23598
x"00",	-- Hex Addr	5C2F	23599
x"00",	-- Hex Addr	5C30	23600
x"00",	-- Hex Addr	5C31	23601
x"00",	-- Hex Addr	5C32	23602
x"00",	-- Hex Addr	5C33	23603
x"00",	-- Hex Addr	5C34	23604
x"00",	-- Hex Addr	5C35	23605
x"00",	-- Hex Addr	5C36	23606
x"00",	-- Hex Addr	5C37	23607
x"00",	-- Hex Addr	5C38	23608
x"00",	-- Hex Addr	5C39	23609
x"00",	-- Hex Addr	5C3A	23610
x"00",	-- Hex Addr	5C3B	23611
x"00",	-- Hex Addr	5C3C	23612
x"00",	-- Hex Addr	5C3D	23613
x"00",	-- Hex Addr	5C3E	23614
x"00",	-- Hex Addr	5C3F	23615
x"00",	-- Hex Addr	5C40	23616
x"00",	-- Hex Addr	5C41	23617
x"00",	-- Hex Addr	5C42	23618
x"00",	-- Hex Addr	5C43	23619
x"00",	-- Hex Addr	5C44	23620
x"00",	-- Hex Addr	5C45	23621
x"00",	-- Hex Addr	5C46	23622
x"00",	-- Hex Addr	5C47	23623
x"00",	-- Hex Addr	5C48	23624
x"00",	-- Hex Addr	5C49	23625
x"00",	-- Hex Addr	5C4A	23626
x"00",	-- Hex Addr	5C4B	23627
x"00",	-- Hex Addr	5C4C	23628
x"00",	-- Hex Addr	5C4D	23629
x"00",	-- Hex Addr	5C4E	23630
x"00",	-- Hex Addr	5C4F	23631
x"00",	-- Hex Addr	5C50	23632
x"00",	-- Hex Addr	5C51	23633
x"00",	-- Hex Addr	5C52	23634
x"00",	-- Hex Addr	5C53	23635
x"00",	-- Hex Addr	5C54	23636
x"00",	-- Hex Addr	5C55	23637
x"00",	-- Hex Addr	5C56	23638
x"00",	-- Hex Addr	5C57	23639
x"00",	-- Hex Addr	5C58	23640
x"00",	-- Hex Addr	5C59	23641
x"00",	-- Hex Addr	5C5A	23642
x"00",	-- Hex Addr	5C5B	23643
x"00",	-- Hex Addr	5C5C	23644
x"00",	-- Hex Addr	5C5D	23645
x"00",	-- Hex Addr	5C5E	23646
x"00",	-- Hex Addr	5C5F	23647
x"00",	-- Hex Addr	5C60	23648
x"00",	-- Hex Addr	5C61	23649
x"00",	-- Hex Addr	5C62	23650
x"00",	-- Hex Addr	5C63	23651
x"00",	-- Hex Addr	5C64	23652
x"00",	-- Hex Addr	5C65	23653
x"00",	-- Hex Addr	5C66	23654
x"00",	-- Hex Addr	5C67	23655
x"00",	-- Hex Addr	5C68	23656
x"00",	-- Hex Addr	5C69	23657
x"00",	-- Hex Addr	5C6A	23658
x"00",	-- Hex Addr	5C6B	23659
x"00",	-- Hex Addr	5C6C	23660
x"00",	-- Hex Addr	5C6D	23661
x"00",	-- Hex Addr	5C6E	23662
x"00",	-- Hex Addr	5C6F	23663
x"00",	-- Hex Addr	5C70	23664
x"00",	-- Hex Addr	5C71	23665
x"00",	-- Hex Addr	5C72	23666
x"00",	-- Hex Addr	5C73	23667
x"00",	-- Hex Addr	5C74	23668
x"00",	-- Hex Addr	5C75	23669
x"00",	-- Hex Addr	5C76	23670
x"00",	-- Hex Addr	5C77	23671
x"00",	-- Hex Addr	5C78	23672
x"00",	-- Hex Addr	5C79	23673
x"00",	-- Hex Addr	5C7A	23674
x"00",	-- Hex Addr	5C7B	23675
x"00",	-- Hex Addr	5C7C	23676
x"00",	-- Hex Addr	5C7D	23677
x"00",	-- Hex Addr	5C7E	23678
x"00",	-- Hex Addr	5C7F	23679
x"00",	-- Hex Addr	5C80	23680
x"00",	-- Hex Addr	5C81	23681
x"00",	-- Hex Addr	5C82	23682
x"00",	-- Hex Addr	5C83	23683
x"00",	-- Hex Addr	5C84	23684
x"00",	-- Hex Addr	5C85	23685
x"00",	-- Hex Addr	5C86	23686
x"00",	-- Hex Addr	5C87	23687
x"00",	-- Hex Addr	5C88	23688
x"00",	-- Hex Addr	5C89	23689
x"00",	-- Hex Addr	5C8A	23690
x"00",	-- Hex Addr	5C8B	23691
x"00",	-- Hex Addr	5C8C	23692
x"00",	-- Hex Addr	5C8D	23693
x"00",	-- Hex Addr	5C8E	23694
x"00",	-- Hex Addr	5C8F	23695
x"00",	-- Hex Addr	5C90	23696
x"00",	-- Hex Addr	5C91	23697
x"00",	-- Hex Addr	5C92	23698
x"00",	-- Hex Addr	5C93	23699
x"00",	-- Hex Addr	5C94	23700
x"00",	-- Hex Addr	5C95	23701
x"00",	-- Hex Addr	5C96	23702
x"00",	-- Hex Addr	5C97	23703
x"00",	-- Hex Addr	5C98	23704
x"00",	-- Hex Addr	5C99	23705
x"00",	-- Hex Addr	5C9A	23706
x"00",	-- Hex Addr	5C9B	23707
x"00",	-- Hex Addr	5C9C	23708
x"00",	-- Hex Addr	5C9D	23709
x"00",	-- Hex Addr	5C9E	23710
x"00",	-- Hex Addr	5C9F	23711
x"00",	-- Hex Addr	5CA0	23712
x"00",	-- Hex Addr	5CA1	23713
x"00",	-- Hex Addr	5CA2	23714
x"00",	-- Hex Addr	5CA3	23715
x"00",	-- Hex Addr	5CA4	23716
x"00",	-- Hex Addr	5CA5	23717
x"00",	-- Hex Addr	5CA6	23718
x"00",	-- Hex Addr	5CA7	23719
x"00",	-- Hex Addr	5CA8	23720
x"00",	-- Hex Addr	5CA9	23721
x"00",	-- Hex Addr	5CAA	23722
x"00",	-- Hex Addr	5CAB	23723
x"00",	-- Hex Addr	5CAC	23724
x"00",	-- Hex Addr	5CAD	23725
x"00",	-- Hex Addr	5CAE	23726
x"00",	-- Hex Addr	5CAF	23727
x"00",	-- Hex Addr	5CB0	23728
x"00",	-- Hex Addr	5CB1	23729
x"00",	-- Hex Addr	5CB2	23730
x"00",	-- Hex Addr	5CB3	23731
x"00",	-- Hex Addr	5CB4	23732
x"00",	-- Hex Addr	5CB5	23733
x"00",	-- Hex Addr	5CB6	23734
x"00",	-- Hex Addr	5CB7	23735
x"00",	-- Hex Addr	5CB8	23736
x"00",	-- Hex Addr	5CB9	23737
x"00",	-- Hex Addr	5CBA	23738
x"00",	-- Hex Addr	5CBB	23739
x"00",	-- Hex Addr	5CBC	23740
x"00",	-- Hex Addr	5CBD	23741
x"00",	-- Hex Addr	5CBE	23742
x"00",	-- Hex Addr	5CBF	23743
x"00",	-- Hex Addr	5CC0	23744
x"00",	-- Hex Addr	5CC1	23745
x"00",	-- Hex Addr	5CC2	23746
x"00",	-- Hex Addr	5CC3	23747
x"00",	-- Hex Addr	5CC4	23748
x"00",	-- Hex Addr	5CC5	23749
x"00",	-- Hex Addr	5CC6	23750
x"00",	-- Hex Addr	5CC7	23751
x"00",	-- Hex Addr	5CC8	23752
x"00",	-- Hex Addr	5CC9	23753
x"00",	-- Hex Addr	5CCA	23754
x"00",	-- Hex Addr	5CCB	23755
x"00",	-- Hex Addr	5CCC	23756
x"00",	-- Hex Addr	5CCD	23757
x"00",	-- Hex Addr	5CCE	23758
x"00",	-- Hex Addr	5CCF	23759
x"00",	-- Hex Addr	5CD0	23760
x"00",	-- Hex Addr	5CD1	23761
x"00",	-- Hex Addr	5CD2	23762
x"00",	-- Hex Addr	5CD3	23763
x"00",	-- Hex Addr	5CD4	23764
x"00",	-- Hex Addr	5CD5	23765
x"00",	-- Hex Addr	5CD6	23766
x"00",	-- Hex Addr	5CD7	23767
x"00",	-- Hex Addr	5CD8	23768
x"00",	-- Hex Addr	5CD9	23769
x"00",	-- Hex Addr	5CDA	23770
x"00",	-- Hex Addr	5CDB	23771
x"00",	-- Hex Addr	5CDC	23772
x"00",	-- Hex Addr	5CDD	23773
x"00",	-- Hex Addr	5CDE	23774
x"00",	-- Hex Addr	5CDF	23775
x"00",	-- Hex Addr	5CE0	23776
x"00",	-- Hex Addr	5CE1	23777
x"00",	-- Hex Addr	5CE2	23778
x"00",	-- Hex Addr	5CE3	23779
x"00",	-- Hex Addr	5CE4	23780
x"00",	-- Hex Addr	5CE5	23781
x"00",	-- Hex Addr	5CE6	23782
x"00",	-- Hex Addr	5CE7	23783
x"00",	-- Hex Addr	5CE8	23784
x"00",	-- Hex Addr	5CE9	23785
x"00",	-- Hex Addr	5CEA	23786
x"00",	-- Hex Addr	5CEB	23787
x"00",	-- Hex Addr	5CEC	23788
x"00",	-- Hex Addr	5CED	23789
x"00",	-- Hex Addr	5CEE	23790
x"00",	-- Hex Addr	5CEF	23791
x"00",	-- Hex Addr	5CF0	23792
x"00",	-- Hex Addr	5CF1	23793
x"00",	-- Hex Addr	5CF2	23794
x"00",	-- Hex Addr	5CF3	23795
x"00",	-- Hex Addr	5CF4	23796
x"00",	-- Hex Addr	5CF5	23797
x"00",	-- Hex Addr	5CF6	23798
x"00",	-- Hex Addr	5CF7	23799
x"00",	-- Hex Addr	5CF8	23800
x"00",	-- Hex Addr	5CF9	23801
x"00",	-- Hex Addr	5CFA	23802
x"00",	-- Hex Addr	5CFB	23803
x"00",	-- Hex Addr	5CFC	23804
x"00",	-- Hex Addr	5CFD	23805
x"00",	-- Hex Addr	5CFE	23806
x"00",	-- Hex Addr	5CFF	23807
x"00",	-- Hex Addr	5D00	23808
x"00",	-- Hex Addr	5D01	23809
x"00",	-- Hex Addr	5D02	23810
x"00",	-- Hex Addr	5D03	23811
x"00",	-- Hex Addr	5D04	23812
x"00",	-- Hex Addr	5D05	23813
x"00",	-- Hex Addr	5D06	23814
x"00",	-- Hex Addr	5D07	23815
x"00",	-- Hex Addr	5D08	23816
x"00",	-- Hex Addr	5D09	23817
x"00",	-- Hex Addr	5D0A	23818
x"00",	-- Hex Addr	5D0B	23819
x"00",	-- Hex Addr	5D0C	23820
x"00",	-- Hex Addr	5D0D	23821
x"00",	-- Hex Addr	5D0E	23822
x"00",	-- Hex Addr	5D0F	23823
x"00",	-- Hex Addr	5D10	23824
x"00",	-- Hex Addr	5D11	23825
x"00",	-- Hex Addr	5D12	23826
x"00",	-- Hex Addr	5D13	23827
x"00",	-- Hex Addr	5D14	23828
x"00",	-- Hex Addr	5D15	23829
x"00",	-- Hex Addr	5D16	23830
x"00",	-- Hex Addr	5D17	23831
x"00",	-- Hex Addr	5D18	23832
x"00",	-- Hex Addr	5D19	23833
x"00",	-- Hex Addr	5D1A	23834
x"00",	-- Hex Addr	5D1B	23835
x"00",	-- Hex Addr	5D1C	23836
x"00",	-- Hex Addr	5D1D	23837
x"00",	-- Hex Addr	5D1E	23838
x"00",	-- Hex Addr	5D1F	23839
x"00",	-- Hex Addr	5D20	23840
x"00",	-- Hex Addr	5D21	23841
x"00",	-- Hex Addr	5D22	23842
x"00",	-- Hex Addr	5D23	23843
x"00",	-- Hex Addr	5D24	23844
x"00",	-- Hex Addr	5D25	23845
x"00",	-- Hex Addr	5D26	23846
x"00",	-- Hex Addr	5D27	23847
x"00",	-- Hex Addr	5D28	23848
x"00",	-- Hex Addr	5D29	23849
x"00",	-- Hex Addr	5D2A	23850
x"00",	-- Hex Addr	5D2B	23851
x"00",	-- Hex Addr	5D2C	23852
x"00",	-- Hex Addr	5D2D	23853
x"00",	-- Hex Addr	5D2E	23854
x"00",	-- Hex Addr	5D2F	23855
x"00",	-- Hex Addr	5D30	23856
x"00",	-- Hex Addr	5D31	23857
x"00",	-- Hex Addr	5D32	23858
x"00",	-- Hex Addr	5D33	23859
x"00",	-- Hex Addr	5D34	23860
x"00",	-- Hex Addr	5D35	23861
x"00",	-- Hex Addr	5D36	23862
x"00",	-- Hex Addr	5D37	23863
x"00",	-- Hex Addr	5D38	23864
x"00",	-- Hex Addr	5D39	23865
x"00",	-- Hex Addr	5D3A	23866
x"00",	-- Hex Addr	5D3B	23867
x"00",	-- Hex Addr	5D3C	23868
x"00",	-- Hex Addr	5D3D	23869
x"00",	-- Hex Addr	5D3E	23870
x"00",	-- Hex Addr	5D3F	23871
x"00",	-- Hex Addr	5D40	23872
x"00",	-- Hex Addr	5D41	23873
x"00",	-- Hex Addr	5D42	23874
x"00",	-- Hex Addr	5D43	23875
x"00",	-- Hex Addr	5D44	23876
x"00",	-- Hex Addr	5D45	23877
x"00",	-- Hex Addr	5D46	23878
x"00",	-- Hex Addr	5D47	23879
x"00",	-- Hex Addr	5D48	23880
x"00",	-- Hex Addr	5D49	23881
x"00",	-- Hex Addr	5D4A	23882
x"00",	-- Hex Addr	5D4B	23883
x"00",	-- Hex Addr	5D4C	23884
x"00",	-- Hex Addr	5D4D	23885
x"00",	-- Hex Addr	5D4E	23886
x"00",	-- Hex Addr	5D4F	23887
x"00",	-- Hex Addr	5D50	23888
x"00",	-- Hex Addr	5D51	23889
x"00",	-- Hex Addr	5D52	23890
x"00",	-- Hex Addr	5D53	23891
x"00",	-- Hex Addr	5D54	23892
x"00",	-- Hex Addr	5D55	23893
x"00",	-- Hex Addr	5D56	23894
x"00",	-- Hex Addr	5D57	23895
x"00",	-- Hex Addr	5D58	23896
x"00",	-- Hex Addr	5D59	23897
x"00",	-- Hex Addr	5D5A	23898
x"00",	-- Hex Addr	5D5B	23899
x"00",	-- Hex Addr	5D5C	23900
x"00",	-- Hex Addr	5D5D	23901
x"00",	-- Hex Addr	5D5E	23902
x"00",	-- Hex Addr	5D5F	23903
x"00",	-- Hex Addr	5D60	23904
x"00",	-- Hex Addr	5D61	23905
x"00",	-- Hex Addr	5D62	23906
x"00",	-- Hex Addr	5D63	23907
x"00",	-- Hex Addr	5D64	23908
x"00",	-- Hex Addr	5D65	23909
x"00",	-- Hex Addr	5D66	23910
x"00",	-- Hex Addr	5D67	23911
x"00",	-- Hex Addr	5D68	23912
x"00",	-- Hex Addr	5D69	23913
x"00",	-- Hex Addr	5D6A	23914
x"00",	-- Hex Addr	5D6B	23915
x"00",	-- Hex Addr	5D6C	23916
x"00",	-- Hex Addr	5D6D	23917
x"00",	-- Hex Addr	5D6E	23918
x"00",	-- Hex Addr	5D6F	23919
x"00",	-- Hex Addr	5D70	23920
x"00",	-- Hex Addr	5D71	23921
x"00",	-- Hex Addr	5D72	23922
x"00",	-- Hex Addr	5D73	23923
x"00",	-- Hex Addr	5D74	23924
x"00",	-- Hex Addr	5D75	23925
x"00",	-- Hex Addr	5D76	23926
x"00",	-- Hex Addr	5D77	23927
x"00",	-- Hex Addr	5D78	23928
x"00",	-- Hex Addr	5D79	23929
x"00",	-- Hex Addr	5D7A	23930
x"00",	-- Hex Addr	5D7B	23931
x"00",	-- Hex Addr	5D7C	23932
x"00",	-- Hex Addr	5D7D	23933
x"00",	-- Hex Addr	5D7E	23934
x"00",	-- Hex Addr	5D7F	23935
x"00",	-- Hex Addr	5D80	23936
x"00",	-- Hex Addr	5D81	23937
x"00",	-- Hex Addr	5D82	23938
x"00",	-- Hex Addr	5D83	23939
x"00",	-- Hex Addr	5D84	23940
x"00",	-- Hex Addr	5D85	23941
x"00",	-- Hex Addr	5D86	23942
x"00",	-- Hex Addr	5D87	23943
x"00",	-- Hex Addr	5D88	23944
x"00",	-- Hex Addr	5D89	23945
x"00",	-- Hex Addr	5D8A	23946
x"00",	-- Hex Addr	5D8B	23947
x"00",	-- Hex Addr	5D8C	23948
x"00",	-- Hex Addr	5D8D	23949
x"00",	-- Hex Addr	5D8E	23950
x"00",	-- Hex Addr	5D8F	23951
x"00",	-- Hex Addr	5D90	23952
x"00",	-- Hex Addr	5D91	23953
x"00",	-- Hex Addr	5D92	23954
x"00",	-- Hex Addr	5D93	23955
x"00",	-- Hex Addr	5D94	23956
x"00",	-- Hex Addr	5D95	23957
x"00",	-- Hex Addr	5D96	23958
x"00",	-- Hex Addr	5D97	23959
x"00",	-- Hex Addr	5D98	23960
x"00",	-- Hex Addr	5D99	23961
x"00",	-- Hex Addr	5D9A	23962
x"00",	-- Hex Addr	5D9B	23963
x"00",	-- Hex Addr	5D9C	23964
x"00",	-- Hex Addr	5D9D	23965
x"00",	-- Hex Addr	5D9E	23966
x"00",	-- Hex Addr	5D9F	23967
x"00",	-- Hex Addr	5DA0	23968
x"00",	-- Hex Addr	5DA1	23969
x"00",	-- Hex Addr	5DA2	23970
x"00",	-- Hex Addr	5DA3	23971
x"00",	-- Hex Addr	5DA4	23972
x"00",	-- Hex Addr	5DA5	23973
x"00",	-- Hex Addr	5DA6	23974
x"00",	-- Hex Addr	5DA7	23975
x"00",	-- Hex Addr	5DA8	23976
x"00",	-- Hex Addr	5DA9	23977
x"00",	-- Hex Addr	5DAA	23978
x"00",	-- Hex Addr	5DAB	23979
x"00",	-- Hex Addr	5DAC	23980
x"00",	-- Hex Addr	5DAD	23981
x"00",	-- Hex Addr	5DAE	23982
x"00",	-- Hex Addr	5DAF	23983
x"00",	-- Hex Addr	5DB0	23984
x"00",	-- Hex Addr	5DB1	23985
x"00",	-- Hex Addr	5DB2	23986
x"00",	-- Hex Addr	5DB3	23987
x"00",	-- Hex Addr	5DB4	23988
x"00",	-- Hex Addr	5DB5	23989
x"00",	-- Hex Addr	5DB6	23990
x"00",	-- Hex Addr	5DB7	23991
x"00",	-- Hex Addr	5DB8	23992
x"00",	-- Hex Addr	5DB9	23993
x"00",	-- Hex Addr	5DBA	23994
x"00",	-- Hex Addr	5DBB	23995
x"00",	-- Hex Addr	5DBC	23996
x"00",	-- Hex Addr	5DBD	23997
x"00",	-- Hex Addr	5DBE	23998
x"00",	-- Hex Addr	5DBF	23999
x"00",	-- Hex Addr	5DC0	24000
x"00",	-- Hex Addr	5DC1	24001
x"00",	-- Hex Addr	5DC2	24002
x"00",	-- Hex Addr	5DC3	24003
x"00",	-- Hex Addr	5DC4	24004
x"00",	-- Hex Addr	5DC5	24005
x"00",	-- Hex Addr	5DC6	24006
x"00",	-- Hex Addr	5DC7	24007
x"00",	-- Hex Addr	5DC8	24008
x"00",	-- Hex Addr	5DC9	24009
x"00",	-- Hex Addr	5DCA	24010
x"00",	-- Hex Addr	5DCB	24011
x"00",	-- Hex Addr	5DCC	24012
x"00",	-- Hex Addr	5DCD	24013
x"00",	-- Hex Addr	5DCE	24014
x"00",	-- Hex Addr	5DCF	24015
x"00",	-- Hex Addr	5DD0	24016
x"00",	-- Hex Addr	5DD1	24017
x"00",	-- Hex Addr	5DD2	24018
x"00",	-- Hex Addr	5DD3	24019
x"00",	-- Hex Addr	5DD4	24020
x"00",	-- Hex Addr	5DD5	24021
x"00",	-- Hex Addr	5DD6	24022
x"00",	-- Hex Addr	5DD7	24023
x"00",	-- Hex Addr	5DD8	24024
x"00",	-- Hex Addr	5DD9	24025
x"00",	-- Hex Addr	5DDA	24026
x"00",	-- Hex Addr	5DDB	24027
x"00",	-- Hex Addr	5DDC	24028
x"00",	-- Hex Addr	5DDD	24029
x"00",	-- Hex Addr	5DDE	24030
x"00",	-- Hex Addr	5DDF	24031
x"00",	-- Hex Addr	5DE0	24032
x"00",	-- Hex Addr	5DE1	24033
x"00",	-- Hex Addr	5DE2	24034
x"00",	-- Hex Addr	5DE3	24035
x"00",	-- Hex Addr	5DE4	24036
x"00",	-- Hex Addr	5DE5	24037
x"00",	-- Hex Addr	5DE6	24038
x"00",	-- Hex Addr	5DE7	24039
x"00",	-- Hex Addr	5DE8	24040
x"00",	-- Hex Addr	5DE9	24041
x"00",	-- Hex Addr	5DEA	24042
x"00",	-- Hex Addr	5DEB	24043
x"00",	-- Hex Addr	5DEC	24044
x"00",	-- Hex Addr	5DED	24045
x"00",	-- Hex Addr	5DEE	24046
x"00",	-- Hex Addr	5DEF	24047
x"00",	-- Hex Addr	5DF0	24048
x"00",	-- Hex Addr	5DF1	24049
x"00",	-- Hex Addr	5DF2	24050
x"00",	-- Hex Addr	5DF3	24051
x"00",	-- Hex Addr	5DF4	24052
x"00",	-- Hex Addr	5DF5	24053
x"00",	-- Hex Addr	5DF6	24054
x"00",	-- Hex Addr	5DF7	24055
x"00",	-- Hex Addr	5DF8	24056
x"00",	-- Hex Addr	5DF9	24057
x"00",	-- Hex Addr	5DFA	24058
x"00",	-- Hex Addr	5DFB	24059
x"00",	-- Hex Addr	5DFC	24060
x"00",	-- Hex Addr	5DFD	24061
x"00",	-- Hex Addr	5DFE	24062
x"00",	-- Hex Addr	5DFF	24063
x"00",	-- Hex Addr	5E00	24064
x"00",	-- Hex Addr	5E01	24065
x"00",	-- Hex Addr	5E02	24066
x"00",	-- Hex Addr	5E03	24067
x"00",	-- Hex Addr	5E04	24068
x"00",	-- Hex Addr	5E05	24069
x"00",	-- Hex Addr	5E06	24070
x"00",	-- Hex Addr	5E07	24071
x"00",	-- Hex Addr	5E08	24072
x"00",	-- Hex Addr	5E09	24073
x"00",	-- Hex Addr	5E0A	24074
x"00",	-- Hex Addr	5E0B	24075
x"00",	-- Hex Addr	5E0C	24076
x"00",	-- Hex Addr	5E0D	24077
x"00",	-- Hex Addr	5E0E	24078
x"00",	-- Hex Addr	5E0F	24079
x"00",	-- Hex Addr	5E10	24080
x"00",	-- Hex Addr	5E11	24081
x"00",	-- Hex Addr	5E12	24082
x"00",	-- Hex Addr	5E13	24083
x"00",	-- Hex Addr	5E14	24084
x"00",	-- Hex Addr	5E15	24085
x"00",	-- Hex Addr	5E16	24086
x"00",	-- Hex Addr	5E17	24087
x"00",	-- Hex Addr	5E18	24088
x"00",	-- Hex Addr	5E19	24089
x"00",	-- Hex Addr	5E1A	24090
x"00",	-- Hex Addr	5E1B	24091
x"00",	-- Hex Addr	5E1C	24092
x"00",	-- Hex Addr	5E1D	24093
x"00",	-- Hex Addr	5E1E	24094
x"00",	-- Hex Addr	5E1F	24095
x"00",	-- Hex Addr	5E20	24096
x"00",	-- Hex Addr	5E21	24097
x"00",	-- Hex Addr	5E22	24098
x"00",	-- Hex Addr	5E23	24099
x"00",	-- Hex Addr	5E24	24100
x"00",	-- Hex Addr	5E25	24101
x"00",	-- Hex Addr	5E26	24102
x"00",	-- Hex Addr	5E27	24103
x"00",	-- Hex Addr	5E28	24104
x"00",	-- Hex Addr	5E29	24105
x"00",	-- Hex Addr	5E2A	24106
x"00",	-- Hex Addr	5E2B	24107
x"00",	-- Hex Addr	5E2C	24108
x"00",	-- Hex Addr	5E2D	24109
x"00",	-- Hex Addr	5E2E	24110
x"00",	-- Hex Addr	5E2F	24111
x"00",	-- Hex Addr	5E30	24112
x"00",	-- Hex Addr	5E31	24113
x"00",	-- Hex Addr	5E32	24114
x"00",	-- Hex Addr	5E33	24115
x"00",	-- Hex Addr	5E34	24116
x"00",	-- Hex Addr	5E35	24117
x"00",	-- Hex Addr	5E36	24118
x"00",	-- Hex Addr	5E37	24119
x"00",	-- Hex Addr	5E38	24120
x"00",	-- Hex Addr	5E39	24121
x"00",	-- Hex Addr	5E3A	24122
x"00",	-- Hex Addr	5E3B	24123
x"00",	-- Hex Addr	5E3C	24124
x"00",	-- Hex Addr	5E3D	24125
x"00",	-- Hex Addr	5E3E	24126
x"00",	-- Hex Addr	5E3F	24127
x"00",	-- Hex Addr	5E40	24128
x"00",	-- Hex Addr	5E41	24129
x"00",	-- Hex Addr	5E42	24130
x"00",	-- Hex Addr	5E43	24131
x"00",	-- Hex Addr	5E44	24132
x"00",	-- Hex Addr	5E45	24133
x"00",	-- Hex Addr	5E46	24134
x"00",	-- Hex Addr	5E47	24135
x"00",	-- Hex Addr	5E48	24136
x"00",	-- Hex Addr	5E49	24137
x"00",	-- Hex Addr	5E4A	24138
x"00",	-- Hex Addr	5E4B	24139
x"00",	-- Hex Addr	5E4C	24140
x"00",	-- Hex Addr	5E4D	24141
x"00",	-- Hex Addr	5E4E	24142
x"00",	-- Hex Addr	5E4F	24143
x"00",	-- Hex Addr	5E50	24144
x"00",	-- Hex Addr	5E51	24145
x"00",	-- Hex Addr	5E52	24146
x"00",	-- Hex Addr	5E53	24147
x"00",	-- Hex Addr	5E54	24148
x"00",	-- Hex Addr	5E55	24149
x"00",	-- Hex Addr	5E56	24150
x"00",	-- Hex Addr	5E57	24151
x"00",	-- Hex Addr	5E58	24152
x"00",	-- Hex Addr	5E59	24153
x"00",	-- Hex Addr	5E5A	24154
x"00",	-- Hex Addr	5E5B	24155
x"00",	-- Hex Addr	5E5C	24156
x"00",	-- Hex Addr	5E5D	24157
x"00",	-- Hex Addr	5E5E	24158
x"00",	-- Hex Addr	5E5F	24159
x"00",	-- Hex Addr	5E60	24160
x"00",	-- Hex Addr	5E61	24161
x"00",	-- Hex Addr	5E62	24162
x"00",	-- Hex Addr	5E63	24163
x"00",	-- Hex Addr	5E64	24164
x"00",	-- Hex Addr	5E65	24165
x"00",	-- Hex Addr	5E66	24166
x"00",	-- Hex Addr	5E67	24167
x"00",	-- Hex Addr	5E68	24168
x"00",	-- Hex Addr	5E69	24169
x"00",	-- Hex Addr	5E6A	24170
x"00",	-- Hex Addr	5E6B	24171
x"00",	-- Hex Addr	5E6C	24172
x"00",	-- Hex Addr	5E6D	24173
x"00",	-- Hex Addr	5E6E	24174
x"00",	-- Hex Addr	5E6F	24175
x"00",	-- Hex Addr	5E70	24176
x"00",	-- Hex Addr	5E71	24177
x"00",	-- Hex Addr	5E72	24178
x"00",	-- Hex Addr	5E73	24179
x"00",	-- Hex Addr	5E74	24180
x"00",	-- Hex Addr	5E75	24181
x"00",	-- Hex Addr	5E76	24182
x"00",	-- Hex Addr	5E77	24183
x"00",	-- Hex Addr	5E78	24184
x"00",	-- Hex Addr	5E79	24185
x"00",	-- Hex Addr	5E7A	24186
x"00",	-- Hex Addr	5E7B	24187
x"00",	-- Hex Addr	5E7C	24188
x"00",	-- Hex Addr	5E7D	24189
x"00",	-- Hex Addr	5E7E	24190
x"00",	-- Hex Addr	5E7F	24191
x"00",	-- Hex Addr	5E80	24192
x"00",	-- Hex Addr	5E81	24193
x"00",	-- Hex Addr	5E82	24194
x"00",	-- Hex Addr	5E83	24195
x"00",	-- Hex Addr	5E84	24196
x"00",	-- Hex Addr	5E85	24197
x"00",	-- Hex Addr	5E86	24198
x"00",	-- Hex Addr	5E87	24199
x"00",	-- Hex Addr	5E88	24200
x"00",	-- Hex Addr	5E89	24201
x"00",	-- Hex Addr	5E8A	24202
x"00",	-- Hex Addr	5E8B	24203
x"00",	-- Hex Addr	5E8C	24204
x"00",	-- Hex Addr	5E8D	24205
x"00",	-- Hex Addr	5E8E	24206
x"00",	-- Hex Addr	5E8F	24207
x"00",	-- Hex Addr	5E90	24208
x"00",	-- Hex Addr	5E91	24209
x"00",	-- Hex Addr	5E92	24210
x"00",	-- Hex Addr	5E93	24211
x"00",	-- Hex Addr	5E94	24212
x"00",	-- Hex Addr	5E95	24213
x"00",	-- Hex Addr	5E96	24214
x"00",	-- Hex Addr	5E97	24215
x"00",	-- Hex Addr	5E98	24216
x"00",	-- Hex Addr	5E99	24217
x"00",	-- Hex Addr	5E9A	24218
x"00",	-- Hex Addr	5E9B	24219
x"00",	-- Hex Addr	5E9C	24220
x"00",	-- Hex Addr	5E9D	24221
x"00",	-- Hex Addr	5E9E	24222
x"00",	-- Hex Addr	5E9F	24223
x"00",	-- Hex Addr	5EA0	24224
x"00",	-- Hex Addr	5EA1	24225
x"00",	-- Hex Addr	5EA2	24226
x"00",	-- Hex Addr	5EA3	24227
x"00",	-- Hex Addr	5EA4	24228
x"00",	-- Hex Addr	5EA5	24229
x"00",	-- Hex Addr	5EA6	24230
x"00",	-- Hex Addr	5EA7	24231
x"00",	-- Hex Addr	5EA8	24232
x"00",	-- Hex Addr	5EA9	24233
x"00",	-- Hex Addr	5EAA	24234
x"00",	-- Hex Addr	5EAB	24235
x"00",	-- Hex Addr	5EAC	24236
x"00",	-- Hex Addr	5EAD	24237
x"00",	-- Hex Addr	5EAE	24238
x"00",	-- Hex Addr	5EAF	24239
x"00",	-- Hex Addr	5EB0	24240
x"00",	-- Hex Addr	5EB1	24241
x"00",	-- Hex Addr	5EB2	24242
x"00",	-- Hex Addr	5EB3	24243
x"00",	-- Hex Addr	5EB4	24244
x"00",	-- Hex Addr	5EB5	24245
x"00",	-- Hex Addr	5EB6	24246
x"00",	-- Hex Addr	5EB7	24247
x"00",	-- Hex Addr	5EB8	24248
x"00",	-- Hex Addr	5EB9	24249
x"00",	-- Hex Addr	5EBA	24250
x"00",	-- Hex Addr	5EBB	24251
x"00",	-- Hex Addr	5EBC	24252
x"00",	-- Hex Addr	5EBD	24253
x"00",	-- Hex Addr	5EBE	24254
x"00",	-- Hex Addr	5EBF	24255
x"00",	-- Hex Addr	5EC0	24256
x"00",	-- Hex Addr	5EC1	24257
x"00",	-- Hex Addr	5EC2	24258
x"00",	-- Hex Addr	5EC3	24259
x"00",	-- Hex Addr	5EC4	24260
x"00",	-- Hex Addr	5EC5	24261
x"00",	-- Hex Addr	5EC6	24262
x"00",	-- Hex Addr	5EC7	24263
x"00",	-- Hex Addr	5EC8	24264
x"00",	-- Hex Addr	5EC9	24265
x"00",	-- Hex Addr	5ECA	24266
x"00",	-- Hex Addr	5ECB	24267
x"00",	-- Hex Addr	5ECC	24268
x"00",	-- Hex Addr	5ECD	24269
x"00",	-- Hex Addr	5ECE	24270
x"00",	-- Hex Addr	5ECF	24271
x"00",	-- Hex Addr	5ED0	24272
x"00",	-- Hex Addr	5ED1	24273
x"00",	-- Hex Addr	5ED2	24274
x"00",	-- Hex Addr	5ED3	24275
x"00",	-- Hex Addr	5ED4	24276
x"00",	-- Hex Addr	5ED5	24277
x"00",	-- Hex Addr	5ED6	24278
x"00",	-- Hex Addr	5ED7	24279
x"00",	-- Hex Addr	5ED8	24280
x"00",	-- Hex Addr	5ED9	24281
x"00",	-- Hex Addr	5EDA	24282
x"00",	-- Hex Addr	5EDB	24283
x"00",	-- Hex Addr	5EDC	24284
x"00",	-- Hex Addr	5EDD	24285
x"00",	-- Hex Addr	5EDE	24286
x"00",	-- Hex Addr	5EDF	24287
x"00",	-- Hex Addr	5EE0	24288
x"00",	-- Hex Addr	5EE1	24289
x"00",	-- Hex Addr	5EE2	24290
x"00",	-- Hex Addr	5EE3	24291
x"00",	-- Hex Addr	5EE4	24292
x"00",	-- Hex Addr	5EE5	24293
x"00",	-- Hex Addr	5EE6	24294
x"00",	-- Hex Addr	5EE7	24295
x"00",	-- Hex Addr	5EE8	24296
x"00",	-- Hex Addr	5EE9	24297
x"00",	-- Hex Addr	5EEA	24298
x"00",	-- Hex Addr	5EEB	24299
x"00",	-- Hex Addr	5EEC	24300
x"00",	-- Hex Addr	5EED	24301
x"00",	-- Hex Addr	5EEE	24302
x"00",	-- Hex Addr	5EEF	24303
x"00",	-- Hex Addr	5EF0	24304
x"00",	-- Hex Addr	5EF1	24305
x"00",	-- Hex Addr	5EF2	24306
x"00",	-- Hex Addr	5EF3	24307
x"00",	-- Hex Addr	5EF4	24308
x"00",	-- Hex Addr	5EF5	24309
x"00",	-- Hex Addr	5EF6	24310
x"00",	-- Hex Addr	5EF7	24311
x"00",	-- Hex Addr	5EF8	24312
x"00",	-- Hex Addr	5EF9	24313
x"00",	-- Hex Addr	5EFA	24314
x"00",	-- Hex Addr	5EFB	24315
x"00",	-- Hex Addr	5EFC	24316
x"00",	-- Hex Addr	5EFD	24317
x"00",	-- Hex Addr	5EFE	24318
x"00",	-- Hex Addr	5EFF	24319
x"00",	-- Hex Addr	5F00	24320
x"00",	-- Hex Addr	5F01	24321
x"00",	-- Hex Addr	5F02	24322
x"00",	-- Hex Addr	5F03	24323
x"00",	-- Hex Addr	5F04	24324
x"00",	-- Hex Addr	5F05	24325
x"00",	-- Hex Addr	5F06	24326
x"00",	-- Hex Addr	5F07	24327
x"00",	-- Hex Addr	5F08	24328
x"00",	-- Hex Addr	5F09	24329
x"00",	-- Hex Addr	5F0A	24330
x"00",	-- Hex Addr	5F0B	24331
x"00",	-- Hex Addr	5F0C	24332
x"00",	-- Hex Addr	5F0D	24333
x"00",	-- Hex Addr	5F0E	24334
x"00",	-- Hex Addr	5F0F	24335
x"00",	-- Hex Addr	5F10	24336
x"00",	-- Hex Addr	5F11	24337
x"00",	-- Hex Addr	5F12	24338
x"00",	-- Hex Addr	5F13	24339
x"00",	-- Hex Addr	5F14	24340
x"00",	-- Hex Addr	5F15	24341
x"00",	-- Hex Addr	5F16	24342
x"00",	-- Hex Addr	5F17	24343
x"00",	-- Hex Addr	5F18	24344
x"00",	-- Hex Addr	5F19	24345
x"00",	-- Hex Addr	5F1A	24346
x"00",	-- Hex Addr	5F1B	24347
x"00",	-- Hex Addr	5F1C	24348
x"00",	-- Hex Addr	5F1D	24349
x"00",	-- Hex Addr	5F1E	24350
x"00",	-- Hex Addr	5F1F	24351
x"00",	-- Hex Addr	5F20	24352
x"00",	-- Hex Addr	5F21	24353
x"00",	-- Hex Addr	5F22	24354
x"00",	-- Hex Addr	5F23	24355
x"00",	-- Hex Addr	5F24	24356
x"00",	-- Hex Addr	5F25	24357
x"00",	-- Hex Addr	5F26	24358
x"00",	-- Hex Addr	5F27	24359
x"00",	-- Hex Addr	5F28	24360
x"00",	-- Hex Addr	5F29	24361
x"00",	-- Hex Addr	5F2A	24362
x"00",	-- Hex Addr	5F2B	24363
x"00",	-- Hex Addr	5F2C	24364
x"00",	-- Hex Addr	5F2D	24365
x"00",	-- Hex Addr	5F2E	24366
x"00",	-- Hex Addr	5F2F	24367
x"00",	-- Hex Addr	5F30	24368
x"00",	-- Hex Addr	5F31	24369
x"00",	-- Hex Addr	5F32	24370
x"00",	-- Hex Addr	5F33	24371
x"00",	-- Hex Addr	5F34	24372
x"00",	-- Hex Addr	5F35	24373
x"00",	-- Hex Addr	5F36	24374
x"00",	-- Hex Addr	5F37	24375
x"00",	-- Hex Addr	5F38	24376
x"00",	-- Hex Addr	5F39	24377
x"00",	-- Hex Addr	5F3A	24378
x"00",	-- Hex Addr	5F3B	24379
x"00",	-- Hex Addr	5F3C	24380
x"00",	-- Hex Addr	5F3D	24381
x"00",	-- Hex Addr	5F3E	24382
x"00",	-- Hex Addr	5F3F	24383
x"00",	-- Hex Addr	5F40	24384
x"00",	-- Hex Addr	5F41	24385
x"00",	-- Hex Addr	5F42	24386
x"00",	-- Hex Addr	5F43	24387
x"00",	-- Hex Addr	5F44	24388
x"00",	-- Hex Addr	5F45	24389
x"00",	-- Hex Addr	5F46	24390
x"00",	-- Hex Addr	5F47	24391
x"00",	-- Hex Addr	5F48	24392
x"00",	-- Hex Addr	5F49	24393
x"00",	-- Hex Addr	5F4A	24394
x"00",	-- Hex Addr	5F4B	24395
x"00",	-- Hex Addr	5F4C	24396
x"00",	-- Hex Addr	5F4D	24397
x"00",	-- Hex Addr	5F4E	24398
x"00",	-- Hex Addr	5F4F	24399
x"00",	-- Hex Addr	5F50	24400
x"00",	-- Hex Addr	5F51	24401
x"00",	-- Hex Addr	5F52	24402
x"00",	-- Hex Addr	5F53	24403
x"00",	-- Hex Addr	5F54	24404
x"00",	-- Hex Addr	5F55	24405
x"00",	-- Hex Addr	5F56	24406
x"00",	-- Hex Addr	5F57	24407
x"00",	-- Hex Addr	5F58	24408
x"00",	-- Hex Addr	5F59	24409
x"00",	-- Hex Addr	5F5A	24410
x"00",	-- Hex Addr	5F5B	24411
x"00",	-- Hex Addr	5F5C	24412
x"00",	-- Hex Addr	5F5D	24413
x"00",	-- Hex Addr	5F5E	24414
x"00",	-- Hex Addr	5F5F	24415
x"00",	-- Hex Addr	5F60	24416
x"00",	-- Hex Addr	5F61	24417
x"00",	-- Hex Addr	5F62	24418
x"00",	-- Hex Addr	5F63	24419
x"00",	-- Hex Addr	5F64	24420
x"00",	-- Hex Addr	5F65	24421
x"00",	-- Hex Addr	5F66	24422
x"00",	-- Hex Addr	5F67	24423
x"00",	-- Hex Addr	5F68	24424
x"00",	-- Hex Addr	5F69	24425
x"00",	-- Hex Addr	5F6A	24426
x"00",	-- Hex Addr	5F6B	24427
x"00",	-- Hex Addr	5F6C	24428
x"00",	-- Hex Addr	5F6D	24429
x"00",	-- Hex Addr	5F6E	24430
x"00",	-- Hex Addr	5F6F	24431
x"00",	-- Hex Addr	5F70	24432
x"00",	-- Hex Addr	5F71	24433
x"00",	-- Hex Addr	5F72	24434
x"00",	-- Hex Addr	5F73	24435
x"00",	-- Hex Addr	5F74	24436
x"00",	-- Hex Addr	5F75	24437
x"00",	-- Hex Addr	5F76	24438
x"00",	-- Hex Addr	5F77	24439
x"00",	-- Hex Addr	5F78	24440
x"00",	-- Hex Addr	5F79	24441
x"00",	-- Hex Addr	5F7A	24442
x"00",	-- Hex Addr	5F7B	24443
x"00",	-- Hex Addr	5F7C	24444
x"00",	-- Hex Addr	5F7D	24445
x"00",	-- Hex Addr	5F7E	24446
x"00",	-- Hex Addr	5F7F	24447
x"00",	-- Hex Addr	5F80	24448
x"00",	-- Hex Addr	5F81	24449
x"00",	-- Hex Addr	5F82	24450
x"00",	-- Hex Addr	5F83	24451
x"00",	-- Hex Addr	5F84	24452
x"00",	-- Hex Addr	5F85	24453
x"00",	-- Hex Addr	5F86	24454
x"00",	-- Hex Addr	5F87	24455
x"00",	-- Hex Addr	5F88	24456
x"00",	-- Hex Addr	5F89	24457
x"00",	-- Hex Addr	5F8A	24458
x"00",	-- Hex Addr	5F8B	24459
x"00",	-- Hex Addr	5F8C	24460
x"00",	-- Hex Addr	5F8D	24461
x"00",	-- Hex Addr	5F8E	24462
x"00",	-- Hex Addr	5F8F	24463
x"00",	-- Hex Addr	5F90	24464
x"00",	-- Hex Addr	5F91	24465
x"00",	-- Hex Addr	5F92	24466
x"00",	-- Hex Addr	5F93	24467
x"00",	-- Hex Addr	5F94	24468
x"00",	-- Hex Addr	5F95	24469
x"00",	-- Hex Addr	5F96	24470
x"00",	-- Hex Addr	5F97	24471
x"00",	-- Hex Addr	5F98	24472
x"00",	-- Hex Addr	5F99	24473
x"00",	-- Hex Addr	5F9A	24474
x"00",	-- Hex Addr	5F9B	24475
x"00",	-- Hex Addr	5F9C	24476
x"00",	-- Hex Addr	5F9D	24477
x"00",	-- Hex Addr	5F9E	24478
x"00",	-- Hex Addr	5F9F	24479
x"00",	-- Hex Addr	5FA0	24480
x"00",	-- Hex Addr	5FA1	24481
x"00",	-- Hex Addr	5FA2	24482
x"00",	-- Hex Addr	5FA3	24483
x"00",	-- Hex Addr	5FA4	24484
x"00",	-- Hex Addr	5FA5	24485
x"00",	-- Hex Addr	5FA6	24486
x"00",	-- Hex Addr	5FA7	24487
x"00",	-- Hex Addr	5FA8	24488
x"00",	-- Hex Addr	5FA9	24489
x"00",	-- Hex Addr	5FAA	24490
x"00",	-- Hex Addr	5FAB	24491
x"00",	-- Hex Addr	5FAC	24492
x"00",	-- Hex Addr	5FAD	24493
x"00",	-- Hex Addr	5FAE	24494
x"00",	-- Hex Addr	5FAF	24495
x"00",	-- Hex Addr	5FB0	24496
x"00",	-- Hex Addr	5FB1	24497
x"00",	-- Hex Addr	5FB2	24498
x"00",	-- Hex Addr	5FB3	24499
x"00",	-- Hex Addr	5FB4	24500
x"00",	-- Hex Addr	5FB5	24501
x"00",	-- Hex Addr	5FB6	24502
x"00",	-- Hex Addr	5FB7	24503
x"00",	-- Hex Addr	5FB8	24504
x"00",	-- Hex Addr	5FB9	24505
x"00",	-- Hex Addr	5FBA	24506
x"00",	-- Hex Addr	5FBB	24507
x"00",	-- Hex Addr	5FBC	24508
x"00",	-- Hex Addr	5FBD	24509
x"00",	-- Hex Addr	5FBE	24510
x"00",	-- Hex Addr	5FBF	24511
x"00",	-- Hex Addr	5FC0	24512
x"00",	-- Hex Addr	5FC1	24513
x"00",	-- Hex Addr	5FC2	24514
x"00",	-- Hex Addr	5FC3	24515
x"00",	-- Hex Addr	5FC4	24516
x"00",	-- Hex Addr	5FC5	24517
x"00",	-- Hex Addr	5FC6	24518
x"00",	-- Hex Addr	5FC7	24519
x"00",	-- Hex Addr	5FC8	24520
x"00",	-- Hex Addr	5FC9	24521
x"00",	-- Hex Addr	5FCA	24522
x"00",	-- Hex Addr	5FCB	24523
x"00",	-- Hex Addr	5FCC	24524
x"00",	-- Hex Addr	5FCD	24525
x"00",	-- Hex Addr	5FCE	24526
x"00",	-- Hex Addr	5FCF	24527
x"00",	-- Hex Addr	5FD0	24528
x"00",	-- Hex Addr	5FD1	24529
x"00",	-- Hex Addr	5FD2	24530
x"00",	-- Hex Addr	5FD3	24531
x"00",	-- Hex Addr	5FD4	24532
x"00",	-- Hex Addr	5FD5	24533
x"00",	-- Hex Addr	5FD6	24534
x"00",	-- Hex Addr	5FD7	24535
x"00",	-- Hex Addr	5FD8	24536
x"00",	-- Hex Addr	5FD9	24537
x"00",	-- Hex Addr	5FDA	24538
x"00",	-- Hex Addr	5FDB	24539
x"00",	-- Hex Addr	5FDC	24540
x"00",	-- Hex Addr	5FDD	24541
x"00",	-- Hex Addr	5FDE	24542
x"00",	-- Hex Addr	5FDF	24543
x"00",	-- Hex Addr	5FE0	24544
x"00",	-- Hex Addr	5FE1	24545
x"00",	-- Hex Addr	5FE2	24546
x"00",	-- Hex Addr	5FE3	24547
x"00",	-- Hex Addr	5FE4	24548
x"00",	-- Hex Addr	5FE5	24549
x"00",	-- Hex Addr	5FE6	24550
x"00",	-- Hex Addr	5FE7	24551
x"00",	-- Hex Addr	5FE8	24552
x"00",	-- Hex Addr	5FE9	24553
x"00",	-- Hex Addr	5FEA	24554
x"00",	-- Hex Addr	5FEB	24555
x"00",	-- Hex Addr	5FEC	24556
x"00",	-- Hex Addr	5FED	24557
x"00",	-- Hex Addr	5FEE	24558
x"00",	-- Hex Addr	5FEF	24559
x"00",	-- Hex Addr	5FF0	24560
x"00",	-- Hex Addr	5FF1	24561
x"00",	-- Hex Addr	5FF2	24562
x"00",	-- Hex Addr	5FF3	24563
x"00",	-- Hex Addr	5FF4	24564
x"00",	-- Hex Addr	5FF5	24565
x"00",	-- Hex Addr	5FF6	24566
x"00",	-- Hex Addr	5FF7	24567
x"00",	-- Hex Addr	5FF8	24568
x"00",	-- Hex Addr	5FF9	24569
x"00",	-- Hex Addr	5FFA	24570
x"00",	-- Hex Addr	5FFB	24571
x"00",	-- Hex Addr	5FFC	24572
x"00",	-- Hex Addr	5FFD	24573
x"00",	-- Hex Addr	5FFE	24574
x"00",	-- Hex Addr	5FFF	24575
x"00",	-- Hex Addr	6000	24576
x"00",	-- Hex Addr	6001	24577
x"00",	-- Hex Addr	6002	24578
x"00",	-- Hex Addr	6003	24579
x"00",	-- Hex Addr	6004	24580
x"00",	-- Hex Addr	6005	24581
x"00",	-- Hex Addr	6006	24582
x"00",	-- Hex Addr	6007	24583
x"00",	-- Hex Addr	6008	24584
x"00",	-- Hex Addr	6009	24585
x"00",	-- Hex Addr	600A	24586
x"00",	-- Hex Addr	600B	24587
x"00",	-- Hex Addr	600C	24588
x"00",	-- Hex Addr	600D	24589
x"00",	-- Hex Addr	600E	24590
x"00",	-- Hex Addr	600F	24591
x"00",	-- Hex Addr	6010	24592
x"00",	-- Hex Addr	6011	24593
x"00",	-- Hex Addr	6012	24594
x"00",	-- Hex Addr	6013	24595
x"00",	-- Hex Addr	6014	24596
x"00",	-- Hex Addr	6015	24597
x"00",	-- Hex Addr	6016	24598
x"00",	-- Hex Addr	6017	24599
x"00",	-- Hex Addr	6018	24600
x"00",	-- Hex Addr	6019	24601
x"00",	-- Hex Addr	601A	24602
x"00",	-- Hex Addr	601B	24603
x"00",	-- Hex Addr	601C	24604
x"00",	-- Hex Addr	601D	24605
x"00",	-- Hex Addr	601E	24606
x"00",	-- Hex Addr	601F	24607
x"00",	-- Hex Addr	6020	24608
x"00",	-- Hex Addr	6021	24609
x"00",	-- Hex Addr	6022	24610
x"00",	-- Hex Addr	6023	24611
x"00",	-- Hex Addr	6024	24612
x"00",	-- Hex Addr	6025	24613
x"00",	-- Hex Addr	6026	24614
x"00",	-- Hex Addr	6027	24615
x"00",	-- Hex Addr	6028	24616
x"00",	-- Hex Addr	6029	24617
x"00",	-- Hex Addr	602A	24618
x"00",	-- Hex Addr	602B	24619
x"00",	-- Hex Addr	602C	24620
x"00",	-- Hex Addr	602D	24621
x"00",	-- Hex Addr	602E	24622
x"00",	-- Hex Addr	602F	24623
x"00",	-- Hex Addr	6030	24624
x"00",	-- Hex Addr	6031	24625
x"00",	-- Hex Addr	6032	24626
x"00",	-- Hex Addr	6033	24627
x"00",	-- Hex Addr	6034	24628
x"00",	-- Hex Addr	6035	24629
x"00",	-- Hex Addr	6036	24630
x"00",	-- Hex Addr	6037	24631
x"00",	-- Hex Addr	6038	24632
x"00",	-- Hex Addr	6039	24633
x"00",	-- Hex Addr	603A	24634
x"00",	-- Hex Addr	603B	24635
x"00",	-- Hex Addr	603C	24636
x"00",	-- Hex Addr	603D	24637
x"00",	-- Hex Addr	603E	24638
x"00",	-- Hex Addr	603F	24639
x"00",	-- Hex Addr	6040	24640
x"00",	-- Hex Addr	6041	24641
x"00",	-- Hex Addr	6042	24642
x"00",	-- Hex Addr	6043	24643
x"00",	-- Hex Addr	6044	24644
x"00",	-- Hex Addr	6045	24645
x"00",	-- Hex Addr	6046	24646
x"00",	-- Hex Addr	6047	24647
x"00",	-- Hex Addr	6048	24648
x"00",	-- Hex Addr	6049	24649
x"00",	-- Hex Addr	604A	24650
x"00",	-- Hex Addr	604B	24651
x"00",	-- Hex Addr	604C	24652
x"00",	-- Hex Addr	604D	24653
x"00",	-- Hex Addr	604E	24654
x"00",	-- Hex Addr	604F	24655
x"00",	-- Hex Addr	6050	24656
x"00",	-- Hex Addr	6051	24657
x"00",	-- Hex Addr	6052	24658
x"00",	-- Hex Addr	6053	24659
x"00",	-- Hex Addr	6054	24660
x"00",	-- Hex Addr	6055	24661
x"00",	-- Hex Addr	6056	24662
x"00",	-- Hex Addr	6057	24663
x"00",	-- Hex Addr	6058	24664
x"00",	-- Hex Addr	6059	24665
x"00",	-- Hex Addr	605A	24666
x"00",	-- Hex Addr	605B	24667
x"00",	-- Hex Addr	605C	24668
x"00",	-- Hex Addr	605D	24669
x"00",	-- Hex Addr	605E	24670
x"00",	-- Hex Addr	605F	24671
x"00",	-- Hex Addr	6060	24672
x"00",	-- Hex Addr	6061	24673
x"00",	-- Hex Addr	6062	24674
x"00",	-- Hex Addr	6063	24675
x"00",	-- Hex Addr	6064	24676
x"00",	-- Hex Addr	6065	24677
x"00",	-- Hex Addr	6066	24678
x"00",	-- Hex Addr	6067	24679
x"00",	-- Hex Addr	6068	24680
x"00",	-- Hex Addr	6069	24681
x"00",	-- Hex Addr	606A	24682
x"00",	-- Hex Addr	606B	24683
x"00",	-- Hex Addr	606C	24684
x"00",	-- Hex Addr	606D	24685
x"00",	-- Hex Addr	606E	24686
x"00",	-- Hex Addr	606F	24687
x"00",	-- Hex Addr	6070	24688
x"00",	-- Hex Addr	6071	24689
x"00",	-- Hex Addr	6072	24690
x"00",	-- Hex Addr	6073	24691
x"00",	-- Hex Addr	6074	24692
x"00",	-- Hex Addr	6075	24693
x"00",	-- Hex Addr	6076	24694
x"00",	-- Hex Addr	6077	24695
x"00",	-- Hex Addr	6078	24696
x"00",	-- Hex Addr	6079	24697
x"00",	-- Hex Addr	607A	24698
x"00",	-- Hex Addr	607B	24699
x"00",	-- Hex Addr	607C	24700
x"00",	-- Hex Addr	607D	24701
x"00",	-- Hex Addr	607E	24702
x"00",	-- Hex Addr	607F	24703
x"00",	-- Hex Addr	6080	24704
x"00",	-- Hex Addr	6081	24705
x"00",	-- Hex Addr	6082	24706
x"00",	-- Hex Addr	6083	24707
x"00",	-- Hex Addr	6084	24708
x"00",	-- Hex Addr	6085	24709
x"00",	-- Hex Addr	6086	24710
x"00",	-- Hex Addr	6087	24711
x"00",	-- Hex Addr	6088	24712
x"00",	-- Hex Addr	6089	24713
x"00",	-- Hex Addr	608A	24714
x"00",	-- Hex Addr	608B	24715
x"00",	-- Hex Addr	608C	24716
x"00",	-- Hex Addr	608D	24717
x"00",	-- Hex Addr	608E	24718
x"00",	-- Hex Addr	608F	24719
x"00",	-- Hex Addr	6090	24720
x"00",	-- Hex Addr	6091	24721
x"00",	-- Hex Addr	6092	24722
x"00",	-- Hex Addr	6093	24723
x"00",	-- Hex Addr	6094	24724
x"00",	-- Hex Addr	6095	24725
x"00",	-- Hex Addr	6096	24726
x"00",	-- Hex Addr	6097	24727
x"00",	-- Hex Addr	6098	24728
x"00",	-- Hex Addr	6099	24729
x"00",	-- Hex Addr	609A	24730
x"00",	-- Hex Addr	609B	24731
x"00",	-- Hex Addr	609C	24732
x"00",	-- Hex Addr	609D	24733
x"00",	-- Hex Addr	609E	24734
x"00",	-- Hex Addr	609F	24735
x"00",	-- Hex Addr	60A0	24736
x"00",	-- Hex Addr	60A1	24737
x"00",	-- Hex Addr	60A2	24738
x"00",	-- Hex Addr	60A3	24739
x"00",	-- Hex Addr	60A4	24740
x"00",	-- Hex Addr	60A5	24741
x"00",	-- Hex Addr	60A6	24742
x"00",	-- Hex Addr	60A7	24743
x"00",	-- Hex Addr	60A8	24744
x"00",	-- Hex Addr	60A9	24745
x"00",	-- Hex Addr	60AA	24746
x"00",	-- Hex Addr	60AB	24747
x"00",	-- Hex Addr	60AC	24748
x"00",	-- Hex Addr	60AD	24749
x"00",	-- Hex Addr	60AE	24750
x"00",	-- Hex Addr	60AF	24751
x"00",	-- Hex Addr	60B0	24752
x"00",	-- Hex Addr	60B1	24753
x"00",	-- Hex Addr	60B2	24754
x"00",	-- Hex Addr	60B3	24755
x"00",	-- Hex Addr	60B4	24756
x"00",	-- Hex Addr	60B5	24757
x"00",	-- Hex Addr	60B6	24758
x"00",	-- Hex Addr	60B7	24759
x"00",	-- Hex Addr	60B8	24760
x"00",	-- Hex Addr	60B9	24761
x"00",	-- Hex Addr	60BA	24762
x"00",	-- Hex Addr	60BB	24763
x"00",	-- Hex Addr	60BC	24764
x"00",	-- Hex Addr	60BD	24765
x"00",	-- Hex Addr	60BE	24766
x"00",	-- Hex Addr	60BF	24767
x"00",	-- Hex Addr	60C0	24768
x"00",	-- Hex Addr	60C1	24769
x"00",	-- Hex Addr	60C2	24770
x"00",	-- Hex Addr	60C3	24771
x"00",	-- Hex Addr	60C4	24772
x"00",	-- Hex Addr	60C5	24773
x"00",	-- Hex Addr	60C6	24774
x"00",	-- Hex Addr	60C7	24775
x"00",	-- Hex Addr	60C8	24776
x"00",	-- Hex Addr	60C9	24777
x"00",	-- Hex Addr	60CA	24778
x"00",	-- Hex Addr	60CB	24779
x"00",	-- Hex Addr	60CC	24780
x"00",	-- Hex Addr	60CD	24781
x"00",	-- Hex Addr	60CE	24782
x"00",	-- Hex Addr	60CF	24783
x"00",	-- Hex Addr	60D0	24784
x"00",	-- Hex Addr	60D1	24785
x"00",	-- Hex Addr	60D2	24786
x"00",	-- Hex Addr	60D3	24787
x"00",	-- Hex Addr	60D4	24788
x"00",	-- Hex Addr	60D5	24789
x"00",	-- Hex Addr	60D6	24790
x"00",	-- Hex Addr	60D7	24791
x"00",	-- Hex Addr	60D8	24792
x"00",	-- Hex Addr	60D9	24793
x"00",	-- Hex Addr	60DA	24794
x"00",	-- Hex Addr	60DB	24795
x"00",	-- Hex Addr	60DC	24796
x"00",	-- Hex Addr	60DD	24797
x"00",	-- Hex Addr	60DE	24798
x"00",	-- Hex Addr	60DF	24799
x"00",	-- Hex Addr	60E0	24800
x"00",	-- Hex Addr	60E1	24801
x"00",	-- Hex Addr	60E2	24802
x"00",	-- Hex Addr	60E3	24803
x"00",	-- Hex Addr	60E4	24804
x"00",	-- Hex Addr	60E5	24805
x"00",	-- Hex Addr	60E6	24806
x"00",	-- Hex Addr	60E7	24807
x"00",	-- Hex Addr	60E8	24808
x"00",	-- Hex Addr	60E9	24809
x"00",	-- Hex Addr	60EA	24810
x"00",	-- Hex Addr	60EB	24811
x"00",	-- Hex Addr	60EC	24812
x"00",	-- Hex Addr	60ED	24813
x"00",	-- Hex Addr	60EE	24814
x"00",	-- Hex Addr	60EF	24815
x"00",	-- Hex Addr	60F0	24816
x"00",	-- Hex Addr	60F1	24817
x"00",	-- Hex Addr	60F2	24818
x"00",	-- Hex Addr	60F3	24819
x"00",	-- Hex Addr	60F4	24820
x"00",	-- Hex Addr	60F5	24821
x"00",	-- Hex Addr	60F6	24822
x"00",	-- Hex Addr	60F7	24823
x"00",	-- Hex Addr	60F8	24824
x"00",	-- Hex Addr	60F9	24825
x"00",	-- Hex Addr	60FA	24826
x"00",	-- Hex Addr	60FB	24827
x"00",	-- Hex Addr	60FC	24828
x"00",	-- Hex Addr	60FD	24829
x"00",	-- Hex Addr	60FE	24830
x"00",	-- Hex Addr	60FF	24831
x"00",	-- Hex Addr	6100	24832
x"00",	-- Hex Addr	6101	24833
x"00",	-- Hex Addr	6102	24834
x"00",	-- Hex Addr	6103	24835
x"00",	-- Hex Addr	6104	24836
x"00",	-- Hex Addr	6105	24837
x"00",	-- Hex Addr	6106	24838
x"00",	-- Hex Addr	6107	24839
x"00",	-- Hex Addr	6108	24840
x"00",	-- Hex Addr	6109	24841
x"00",	-- Hex Addr	610A	24842
x"00",	-- Hex Addr	610B	24843
x"00",	-- Hex Addr	610C	24844
x"00",	-- Hex Addr	610D	24845
x"00",	-- Hex Addr	610E	24846
x"00",	-- Hex Addr	610F	24847
x"00",	-- Hex Addr	6110	24848
x"00",	-- Hex Addr	6111	24849
x"00",	-- Hex Addr	6112	24850
x"00",	-- Hex Addr	6113	24851
x"00",	-- Hex Addr	6114	24852
x"00",	-- Hex Addr	6115	24853
x"00",	-- Hex Addr	6116	24854
x"00",	-- Hex Addr	6117	24855
x"00",	-- Hex Addr	6118	24856
x"00",	-- Hex Addr	6119	24857
x"00",	-- Hex Addr	611A	24858
x"00",	-- Hex Addr	611B	24859
x"00",	-- Hex Addr	611C	24860
x"00",	-- Hex Addr	611D	24861
x"00",	-- Hex Addr	611E	24862
x"00",	-- Hex Addr	611F	24863
x"00",	-- Hex Addr	6120	24864
x"00",	-- Hex Addr	6121	24865
x"00",	-- Hex Addr	6122	24866
x"00",	-- Hex Addr	6123	24867
x"00",	-- Hex Addr	6124	24868
x"00",	-- Hex Addr	6125	24869
x"00",	-- Hex Addr	6126	24870
x"00",	-- Hex Addr	6127	24871
x"00",	-- Hex Addr	6128	24872
x"00",	-- Hex Addr	6129	24873
x"00",	-- Hex Addr	612A	24874
x"00",	-- Hex Addr	612B	24875
x"00",	-- Hex Addr	612C	24876
x"00",	-- Hex Addr	612D	24877
x"00",	-- Hex Addr	612E	24878
x"00",	-- Hex Addr	612F	24879
x"00",	-- Hex Addr	6130	24880
x"00",	-- Hex Addr	6131	24881
x"00",	-- Hex Addr	6132	24882
x"00",	-- Hex Addr	6133	24883
x"00",	-- Hex Addr	6134	24884
x"00",	-- Hex Addr	6135	24885
x"00",	-- Hex Addr	6136	24886
x"00",	-- Hex Addr	6137	24887
x"00",	-- Hex Addr	6138	24888
x"00",	-- Hex Addr	6139	24889
x"00",	-- Hex Addr	613A	24890
x"00",	-- Hex Addr	613B	24891
x"00",	-- Hex Addr	613C	24892
x"00",	-- Hex Addr	613D	24893
x"00",	-- Hex Addr	613E	24894
x"00",	-- Hex Addr	613F	24895
x"00",	-- Hex Addr	6140	24896
x"00",	-- Hex Addr	6141	24897
x"00",	-- Hex Addr	6142	24898
x"00",	-- Hex Addr	6143	24899
x"00",	-- Hex Addr	6144	24900
x"00",	-- Hex Addr	6145	24901
x"00",	-- Hex Addr	6146	24902
x"00",	-- Hex Addr	6147	24903
x"00",	-- Hex Addr	6148	24904
x"00",	-- Hex Addr	6149	24905
x"00",	-- Hex Addr	614A	24906
x"00",	-- Hex Addr	614B	24907
x"00",	-- Hex Addr	614C	24908
x"00",	-- Hex Addr	614D	24909
x"00",	-- Hex Addr	614E	24910
x"00",	-- Hex Addr	614F	24911
x"00",	-- Hex Addr	6150	24912
x"00",	-- Hex Addr	6151	24913
x"00",	-- Hex Addr	6152	24914
x"00",	-- Hex Addr	6153	24915
x"00",	-- Hex Addr	6154	24916
x"00",	-- Hex Addr	6155	24917
x"00",	-- Hex Addr	6156	24918
x"00",	-- Hex Addr	6157	24919
x"00",	-- Hex Addr	6158	24920
x"00",	-- Hex Addr	6159	24921
x"00",	-- Hex Addr	615A	24922
x"00",	-- Hex Addr	615B	24923
x"00",	-- Hex Addr	615C	24924
x"00",	-- Hex Addr	615D	24925
x"00",	-- Hex Addr	615E	24926
x"00",	-- Hex Addr	615F	24927
x"00",	-- Hex Addr	6160	24928
x"00",	-- Hex Addr	6161	24929
x"00",	-- Hex Addr	6162	24930
x"00",	-- Hex Addr	6163	24931
x"00",	-- Hex Addr	6164	24932
x"00",	-- Hex Addr	6165	24933
x"00",	-- Hex Addr	6166	24934
x"00",	-- Hex Addr	6167	24935
x"00",	-- Hex Addr	6168	24936
x"00",	-- Hex Addr	6169	24937
x"00",	-- Hex Addr	616A	24938
x"00",	-- Hex Addr	616B	24939
x"00",	-- Hex Addr	616C	24940
x"00",	-- Hex Addr	616D	24941
x"00",	-- Hex Addr	616E	24942
x"00",	-- Hex Addr	616F	24943
x"00",	-- Hex Addr	6170	24944
x"00",	-- Hex Addr	6171	24945
x"00",	-- Hex Addr	6172	24946
x"00",	-- Hex Addr	6173	24947
x"00",	-- Hex Addr	6174	24948
x"00",	-- Hex Addr	6175	24949
x"00",	-- Hex Addr	6176	24950
x"00",	-- Hex Addr	6177	24951
x"00",	-- Hex Addr	6178	24952
x"00",	-- Hex Addr	6179	24953
x"00",	-- Hex Addr	617A	24954
x"00",	-- Hex Addr	617B	24955
x"00",	-- Hex Addr	617C	24956
x"00",	-- Hex Addr	617D	24957
x"00",	-- Hex Addr	617E	24958
x"00",	-- Hex Addr	617F	24959
x"00",	-- Hex Addr	6180	24960
x"00",	-- Hex Addr	6181	24961
x"00",	-- Hex Addr	6182	24962
x"00",	-- Hex Addr	6183	24963
x"00",	-- Hex Addr	6184	24964
x"00",	-- Hex Addr	6185	24965
x"00",	-- Hex Addr	6186	24966
x"00",	-- Hex Addr	6187	24967
x"00",	-- Hex Addr	6188	24968
x"00",	-- Hex Addr	6189	24969
x"00",	-- Hex Addr	618A	24970
x"00",	-- Hex Addr	618B	24971
x"00",	-- Hex Addr	618C	24972
x"00",	-- Hex Addr	618D	24973
x"00",	-- Hex Addr	618E	24974
x"00",	-- Hex Addr	618F	24975
x"00",	-- Hex Addr	6190	24976
x"00",	-- Hex Addr	6191	24977
x"00",	-- Hex Addr	6192	24978
x"00",	-- Hex Addr	6193	24979
x"00",	-- Hex Addr	6194	24980
x"00",	-- Hex Addr	6195	24981
x"00",	-- Hex Addr	6196	24982
x"00",	-- Hex Addr	6197	24983
x"00",	-- Hex Addr	6198	24984
x"00",	-- Hex Addr	6199	24985
x"00",	-- Hex Addr	619A	24986
x"00",	-- Hex Addr	619B	24987
x"00",	-- Hex Addr	619C	24988
x"00",	-- Hex Addr	619D	24989
x"00",	-- Hex Addr	619E	24990
x"00",	-- Hex Addr	619F	24991
x"00",	-- Hex Addr	61A0	24992
x"00",	-- Hex Addr	61A1	24993
x"00",	-- Hex Addr	61A2	24994
x"00",	-- Hex Addr	61A3	24995
x"00",	-- Hex Addr	61A4	24996
x"00",	-- Hex Addr	61A5	24997
x"00",	-- Hex Addr	61A6	24998
x"00",	-- Hex Addr	61A7	24999
x"00",	-- Hex Addr	61A8	25000
x"00",	-- Hex Addr	61A9	25001
x"00",	-- Hex Addr	61AA	25002
x"00",	-- Hex Addr	61AB	25003
x"00",	-- Hex Addr	61AC	25004
x"00",	-- Hex Addr	61AD	25005
x"00",	-- Hex Addr	61AE	25006
x"00",	-- Hex Addr	61AF	25007
x"00",	-- Hex Addr	61B0	25008
x"00",	-- Hex Addr	61B1	25009
x"00",	-- Hex Addr	61B2	25010
x"00",	-- Hex Addr	61B3	25011
x"00",	-- Hex Addr	61B4	25012
x"00",	-- Hex Addr	61B5	25013
x"00",	-- Hex Addr	61B6	25014
x"00",	-- Hex Addr	61B7	25015
x"00",	-- Hex Addr	61B8	25016
x"00",	-- Hex Addr	61B9	25017
x"00",	-- Hex Addr	61BA	25018
x"00",	-- Hex Addr	61BB	25019
x"00",	-- Hex Addr	61BC	25020
x"00",	-- Hex Addr	61BD	25021
x"00",	-- Hex Addr	61BE	25022
x"00",	-- Hex Addr	61BF	25023
x"00",	-- Hex Addr	61C0	25024
x"00",	-- Hex Addr	61C1	25025
x"00",	-- Hex Addr	61C2	25026
x"00",	-- Hex Addr	61C3	25027
x"00",	-- Hex Addr	61C4	25028
x"00",	-- Hex Addr	61C5	25029
x"00",	-- Hex Addr	61C6	25030
x"00",	-- Hex Addr	61C7	25031
x"00",	-- Hex Addr	61C8	25032
x"00",	-- Hex Addr	61C9	25033
x"00",	-- Hex Addr	61CA	25034
x"00",	-- Hex Addr	61CB	25035
x"00",	-- Hex Addr	61CC	25036
x"00",	-- Hex Addr	61CD	25037
x"00",	-- Hex Addr	61CE	25038
x"00",	-- Hex Addr	61CF	25039
x"00",	-- Hex Addr	61D0	25040
x"00",	-- Hex Addr	61D1	25041
x"00",	-- Hex Addr	61D2	25042
x"00",	-- Hex Addr	61D3	25043
x"00",	-- Hex Addr	61D4	25044
x"00",	-- Hex Addr	61D5	25045
x"00",	-- Hex Addr	61D6	25046
x"00",	-- Hex Addr	61D7	25047
x"00",	-- Hex Addr	61D8	25048
x"00",	-- Hex Addr	61D9	25049
x"00",	-- Hex Addr	61DA	25050
x"00",	-- Hex Addr	61DB	25051
x"00",	-- Hex Addr	61DC	25052
x"00",	-- Hex Addr	61DD	25053
x"00",	-- Hex Addr	61DE	25054
x"00",	-- Hex Addr	61DF	25055
x"00",	-- Hex Addr	61E0	25056
x"00",	-- Hex Addr	61E1	25057
x"00",	-- Hex Addr	61E2	25058
x"00",	-- Hex Addr	61E3	25059
x"00",	-- Hex Addr	61E4	25060
x"00",	-- Hex Addr	61E5	25061
x"00",	-- Hex Addr	61E6	25062
x"00",	-- Hex Addr	61E7	25063
x"00",	-- Hex Addr	61E8	25064
x"00",	-- Hex Addr	61E9	25065
x"00",	-- Hex Addr	61EA	25066
x"00",	-- Hex Addr	61EB	25067
x"00",	-- Hex Addr	61EC	25068
x"00",	-- Hex Addr	61ED	25069
x"00",	-- Hex Addr	61EE	25070
x"00",	-- Hex Addr	61EF	25071
x"00",	-- Hex Addr	61F0	25072
x"00",	-- Hex Addr	61F1	25073
x"00",	-- Hex Addr	61F2	25074
x"00",	-- Hex Addr	61F3	25075
x"00",	-- Hex Addr	61F4	25076
x"00",	-- Hex Addr	61F5	25077
x"00",	-- Hex Addr	61F6	25078
x"00",	-- Hex Addr	61F7	25079
x"00",	-- Hex Addr	61F8	25080
x"00",	-- Hex Addr	61F9	25081
x"00",	-- Hex Addr	61FA	25082
x"00",	-- Hex Addr	61FB	25083
x"00",	-- Hex Addr	61FC	25084
x"00",	-- Hex Addr	61FD	25085
x"00",	-- Hex Addr	61FE	25086
x"00",	-- Hex Addr	61FF	25087
x"00",	-- Hex Addr	6200	25088
x"00",	-- Hex Addr	6201	25089
x"00",	-- Hex Addr	6202	25090
x"00",	-- Hex Addr	6203	25091
x"00",	-- Hex Addr	6204	25092
x"00",	-- Hex Addr	6205	25093
x"00",	-- Hex Addr	6206	25094
x"00",	-- Hex Addr	6207	25095
x"00",	-- Hex Addr	6208	25096
x"00",	-- Hex Addr	6209	25097
x"00",	-- Hex Addr	620A	25098
x"00",	-- Hex Addr	620B	25099
x"00",	-- Hex Addr	620C	25100
x"00",	-- Hex Addr	620D	25101
x"00",	-- Hex Addr	620E	25102
x"00",	-- Hex Addr	620F	25103
x"00",	-- Hex Addr	6210	25104
x"00",	-- Hex Addr	6211	25105
x"00",	-- Hex Addr	6212	25106
x"00",	-- Hex Addr	6213	25107
x"00",	-- Hex Addr	6214	25108
x"00",	-- Hex Addr	6215	25109
x"00",	-- Hex Addr	6216	25110
x"00",	-- Hex Addr	6217	25111
x"00",	-- Hex Addr	6218	25112
x"00",	-- Hex Addr	6219	25113
x"00",	-- Hex Addr	621A	25114
x"00",	-- Hex Addr	621B	25115
x"00",	-- Hex Addr	621C	25116
x"00",	-- Hex Addr	621D	25117
x"00",	-- Hex Addr	621E	25118
x"00",	-- Hex Addr	621F	25119
x"00",	-- Hex Addr	6220	25120
x"00",	-- Hex Addr	6221	25121
x"00",	-- Hex Addr	6222	25122
x"00",	-- Hex Addr	6223	25123
x"00",	-- Hex Addr	6224	25124
x"00",	-- Hex Addr	6225	25125
x"00",	-- Hex Addr	6226	25126
x"00",	-- Hex Addr	6227	25127
x"00",	-- Hex Addr	6228	25128
x"00",	-- Hex Addr	6229	25129
x"00",	-- Hex Addr	622A	25130
x"00",	-- Hex Addr	622B	25131
x"00",	-- Hex Addr	622C	25132
x"00",	-- Hex Addr	622D	25133
x"00",	-- Hex Addr	622E	25134
x"00",	-- Hex Addr	622F	25135
x"00",	-- Hex Addr	6230	25136
x"00",	-- Hex Addr	6231	25137
x"00",	-- Hex Addr	6232	25138
x"00",	-- Hex Addr	6233	25139
x"00",	-- Hex Addr	6234	25140
x"00",	-- Hex Addr	6235	25141
x"00",	-- Hex Addr	6236	25142
x"00",	-- Hex Addr	6237	25143
x"00",	-- Hex Addr	6238	25144
x"00",	-- Hex Addr	6239	25145
x"00",	-- Hex Addr	623A	25146
x"00",	-- Hex Addr	623B	25147
x"00",	-- Hex Addr	623C	25148
x"00",	-- Hex Addr	623D	25149
x"00",	-- Hex Addr	623E	25150
x"00",	-- Hex Addr	623F	25151
x"00",	-- Hex Addr	6240	25152
x"00",	-- Hex Addr	6241	25153
x"00",	-- Hex Addr	6242	25154
x"00",	-- Hex Addr	6243	25155
x"00",	-- Hex Addr	6244	25156
x"00",	-- Hex Addr	6245	25157
x"00",	-- Hex Addr	6246	25158
x"00",	-- Hex Addr	6247	25159
x"00",	-- Hex Addr	6248	25160
x"00",	-- Hex Addr	6249	25161
x"00",	-- Hex Addr	624A	25162
x"00",	-- Hex Addr	624B	25163
x"00",	-- Hex Addr	624C	25164
x"00",	-- Hex Addr	624D	25165
x"00",	-- Hex Addr	624E	25166
x"00",	-- Hex Addr	624F	25167
x"00",	-- Hex Addr	6250	25168
x"00",	-- Hex Addr	6251	25169
x"00",	-- Hex Addr	6252	25170
x"00",	-- Hex Addr	6253	25171
x"00",	-- Hex Addr	6254	25172
x"00",	-- Hex Addr	6255	25173
x"00",	-- Hex Addr	6256	25174
x"00",	-- Hex Addr	6257	25175
x"00",	-- Hex Addr	6258	25176
x"00",	-- Hex Addr	6259	25177
x"00",	-- Hex Addr	625A	25178
x"00",	-- Hex Addr	625B	25179
x"00",	-- Hex Addr	625C	25180
x"00",	-- Hex Addr	625D	25181
x"00",	-- Hex Addr	625E	25182
x"00",	-- Hex Addr	625F	25183
x"00",	-- Hex Addr	6260	25184
x"00",	-- Hex Addr	6261	25185
x"00",	-- Hex Addr	6262	25186
x"00",	-- Hex Addr	6263	25187
x"00",	-- Hex Addr	6264	25188
x"00",	-- Hex Addr	6265	25189
x"00",	-- Hex Addr	6266	25190
x"00",	-- Hex Addr	6267	25191
x"00",	-- Hex Addr	6268	25192
x"00",	-- Hex Addr	6269	25193
x"00",	-- Hex Addr	626A	25194
x"00",	-- Hex Addr	626B	25195
x"00",	-- Hex Addr	626C	25196
x"00",	-- Hex Addr	626D	25197
x"00",	-- Hex Addr	626E	25198
x"00",	-- Hex Addr	626F	25199
x"00",	-- Hex Addr	6270	25200
x"00",	-- Hex Addr	6271	25201
x"00",	-- Hex Addr	6272	25202
x"00",	-- Hex Addr	6273	25203
x"00",	-- Hex Addr	6274	25204
x"00",	-- Hex Addr	6275	25205
x"00",	-- Hex Addr	6276	25206
x"00",	-- Hex Addr	6277	25207
x"00",	-- Hex Addr	6278	25208
x"00",	-- Hex Addr	6279	25209
x"00",	-- Hex Addr	627A	25210
x"00",	-- Hex Addr	627B	25211
x"00",	-- Hex Addr	627C	25212
x"00",	-- Hex Addr	627D	25213
x"00",	-- Hex Addr	627E	25214
x"00",	-- Hex Addr	627F	25215
x"00",	-- Hex Addr	6280	25216
x"00",	-- Hex Addr	6281	25217
x"00",	-- Hex Addr	6282	25218
x"00",	-- Hex Addr	6283	25219
x"00",	-- Hex Addr	6284	25220
x"00",	-- Hex Addr	6285	25221
x"00",	-- Hex Addr	6286	25222
x"00",	-- Hex Addr	6287	25223
x"00",	-- Hex Addr	6288	25224
x"00",	-- Hex Addr	6289	25225
x"00",	-- Hex Addr	628A	25226
x"00",	-- Hex Addr	628B	25227
x"00",	-- Hex Addr	628C	25228
x"00",	-- Hex Addr	628D	25229
x"00",	-- Hex Addr	628E	25230
x"00",	-- Hex Addr	628F	25231
x"00",	-- Hex Addr	6290	25232
x"00",	-- Hex Addr	6291	25233
x"00",	-- Hex Addr	6292	25234
x"00",	-- Hex Addr	6293	25235
x"00",	-- Hex Addr	6294	25236
x"00",	-- Hex Addr	6295	25237
x"00",	-- Hex Addr	6296	25238
x"00",	-- Hex Addr	6297	25239
x"00",	-- Hex Addr	6298	25240
x"00",	-- Hex Addr	6299	25241
x"00",	-- Hex Addr	629A	25242
x"00",	-- Hex Addr	629B	25243
x"00",	-- Hex Addr	629C	25244
x"00",	-- Hex Addr	629D	25245
x"00",	-- Hex Addr	629E	25246
x"00",	-- Hex Addr	629F	25247
x"00",	-- Hex Addr	62A0	25248
x"00",	-- Hex Addr	62A1	25249
x"00",	-- Hex Addr	62A2	25250
x"00",	-- Hex Addr	62A3	25251
x"00",	-- Hex Addr	62A4	25252
x"00",	-- Hex Addr	62A5	25253
x"00",	-- Hex Addr	62A6	25254
x"00",	-- Hex Addr	62A7	25255
x"00",	-- Hex Addr	62A8	25256
x"00",	-- Hex Addr	62A9	25257
x"00",	-- Hex Addr	62AA	25258
x"00",	-- Hex Addr	62AB	25259
x"00",	-- Hex Addr	62AC	25260
x"00",	-- Hex Addr	62AD	25261
x"00",	-- Hex Addr	62AE	25262
x"00",	-- Hex Addr	62AF	25263
x"00",	-- Hex Addr	62B0	25264
x"00",	-- Hex Addr	62B1	25265
x"00",	-- Hex Addr	62B2	25266
x"00",	-- Hex Addr	62B3	25267
x"00",	-- Hex Addr	62B4	25268
x"00",	-- Hex Addr	62B5	25269
x"00",	-- Hex Addr	62B6	25270
x"00",	-- Hex Addr	62B7	25271
x"00",	-- Hex Addr	62B8	25272
x"00",	-- Hex Addr	62B9	25273
x"00",	-- Hex Addr	62BA	25274
x"00",	-- Hex Addr	62BB	25275
x"00",	-- Hex Addr	62BC	25276
x"00",	-- Hex Addr	62BD	25277
x"00",	-- Hex Addr	62BE	25278
x"00",	-- Hex Addr	62BF	25279
x"00",	-- Hex Addr	62C0	25280
x"00",	-- Hex Addr	62C1	25281
x"00",	-- Hex Addr	62C2	25282
x"00",	-- Hex Addr	62C3	25283
x"00",	-- Hex Addr	62C4	25284
x"00",	-- Hex Addr	62C5	25285
x"00",	-- Hex Addr	62C6	25286
x"00",	-- Hex Addr	62C7	25287
x"00",	-- Hex Addr	62C8	25288
x"00",	-- Hex Addr	62C9	25289
x"00",	-- Hex Addr	62CA	25290
x"00",	-- Hex Addr	62CB	25291
x"00",	-- Hex Addr	62CC	25292
x"00",	-- Hex Addr	62CD	25293
x"00",	-- Hex Addr	62CE	25294
x"00",	-- Hex Addr	62CF	25295
x"00",	-- Hex Addr	62D0	25296
x"00",	-- Hex Addr	62D1	25297
x"00",	-- Hex Addr	62D2	25298
x"00",	-- Hex Addr	62D3	25299
x"00",	-- Hex Addr	62D4	25300
x"00",	-- Hex Addr	62D5	25301
x"00",	-- Hex Addr	62D6	25302
x"00",	-- Hex Addr	62D7	25303
x"00",	-- Hex Addr	62D8	25304
x"00",	-- Hex Addr	62D9	25305
x"00",	-- Hex Addr	62DA	25306
x"00",	-- Hex Addr	62DB	25307
x"00",	-- Hex Addr	62DC	25308
x"00",	-- Hex Addr	62DD	25309
x"00",	-- Hex Addr	62DE	25310
x"00",	-- Hex Addr	62DF	25311
x"00",	-- Hex Addr	62E0	25312
x"00",	-- Hex Addr	62E1	25313
x"00",	-- Hex Addr	62E2	25314
x"00",	-- Hex Addr	62E3	25315
x"00",	-- Hex Addr	62E4	25316
x"00",	-- Hex Addr	62E5	25317
x"00",	-- Hex Addr	62E6	25318
x"00",	-- Hex Addr	62E7	25319
x"00",	-- Hex Addr	62E8	25320
x"00",	-- Hex Addr	62E9	25321
x"00",	-- Hex Addr	62EA	25322
x"00",	-- Hex Addr	62EB	25323
x"00",	-- Hex Addr	62EC	25324
x"00",	-- Hex Addr	62ED	25325
x"00",	-- Hex Addr	62EE	25326
x"00",	-- Hex Addr	62EF	25327
x"00",	-- Hex Addr	62F0	25328
x"00",	-- Hex Addr	62F1	25329
x"00",	-- Hex Addr	62F2	25330
x"00",	-- Hex Addr	62F3	25331
x"00",	-- Hex Addr	62F4	25332
x"00",	-- Hex Addr	62F5	25333
x"00",	-- Hex Addr	62F6	25334
x"00",	-- Hex Addr	62F7	25335
x"00",	-- Hex Addr	62F8	25336
x"00",	-- Hex Addr	62F9	25337
x"00",	-- Hex Addr	62FA	25338
x"00",	-- Hex Addr	62FB	25339
x"00",	-- Hex Addr	62FC	25340
x"00",	-- Hex Addr	62FD	25341
x"00",	-- Hex Addr	62FE	25342
x"00",	-- Hex Addr	62FF	25343
x"00",	-- Hex Addr	6300	25344
x"00",	-- Hex Addr	6301	25345
x"00",	-- Hex Addr	6302	25346
x"00",	-- Hex Addr	6303	25347
x"00",	-- Hex Addr	6304	25348
x"00",	-- Hex Addr	6305	25349
x"00",	-- Hex Addr	6306	25350
x"00",	-- Hex Addr	6307	25351
x"00",	-- Hex Addr	6308	25352
x"00",	-- Hex Addr	6309	25353
x"00",	-- Hex Addr	630A	25354
x"00",	-- Hex Addr	630B	25355
x"00",	-- Hex Addr	630C	25356
x"00",	-- Hex Addr	630D	25357
x"00",	-- Hex Addr	630E	25358
x"00",	-- Hex Addr	630F	25359
x"00",	-- Hex Addr	6310	25360
x"00",	-- Hex Addr	6311	25361
x"00",	-- Hex Addr	6312	25362
x"00",	-- Hex Addr	6313	25363
x"00",	-- Hex Addr	6314	25364
x"00",	-- Hex Addr	6315	25365
x"00",	-- Hex Addr	6316	25366
x"00",	-- Hex Addr	6317	25367
x"00",	-- Hex Addr	6318	25368
x"00",	-- Hex Addr	6319	25369
x"00",	-- Hex Addr	631A	25370
x"00",	-- Hex Addr	631B	25371
x"00",	-- Hex Addr	631C	25372
x"00",	-- Hex Addr	631D	25373
x"00",	-- Hex Addr	631E	25374
x"00",	-- Hex Addr	631F	25375
x"00",	-- Hex Addr	6320	25376
x"00",	-- Hex Addr	6321	25377
x"00",	-- Hex Addr	6322	25378
x"00",	-- Hex Addr	6323	25379
x"00",	-- Hex Addr	6324	25380
x"00",	-- Hex Addr	6325	25381
x"00",	-- Hex Addr	6326	25382
x"00",	-- Hex Addr	6327	25383
x"00",	-- Hex Addr	6328	25384
x"00",	-- Hex Addr	6329	25385
x"00",	-- Hex Addr	632A	25386
x"00",	-- Hex Addr	632B	25387
x"00",	-- Hex Addr	632C	25388
x"00",	-- Hex Addr	632D	25389
x"00",	-- Hex Addr	632E	25390
x"00",	-- Hex Addr	632F	25391
x"00",	-- Hex Addr	6330	25392
x"00",	-- Hex Addr	6331	25393
x"00",	-- Hex Addr	6332	25394
x"00",	-- Hex Addr	6333	25395
x"00",	-- Hex Addr	6334	25396
x"00",	-- Hex Addr	6335	25397
x"00",	-- Hex Addr	6336	25398
x"00",	-- Hex Addr	6337	25399
x"00",	-- Hex Addr	6338	25400
x"00",	-- Hex Addr	6339	25401
x"00",	-- Hex Addr	633A	25402
x"00",	-- Hex Addr	633B	25403
x"00",	-- Hex Addr	633C	25404
x"00",	-- Hex Addr	633D	25405
x"00",	-- Hex Addr	633E	25406
x"00",	-- Hex Addr	633F	25407
x"00",	-- Hex Addr	6340	25408
x"00",	-- Hex Addr	6341	25409
x"00",	-- Hex Addr	6342	25410
x"00",	-- Hex Addr	6343	25411
x"00",	-- Hex Addr	6344	25412
x"00",	-- Hex Addr	6345	25413
x"00",	-- Hex Addr	6346	25414
x"00",	-- Hex Addr	6347	25415
x"00",	-- Hex Addr	6348	25416
x"00",	-- Hex Addr	6349	25417
x"00",	-- Hex Addr	634A	25418
x"00",	-- Hex Addr	634B	25419
x"00",	-- Hex Addr	634C	25420
x"00",	-- Hex Addr	634D	25421
x"00",	-- Hex Addr	634E	25422
x"00",	-- Hex Addr	634F	25423
x"00",	-- Hex Addr	6350	25424
x"00",	-- Hex Addr	6351	25425
x"00",	-- Hex Addr	6352	25426
x"00",	-- Hex Addr	6353	25427
x"00",	-- Hex Addr	6354	25428
x"00",	-- Hex Addr	6355	25429
x"00",	-- Hex Addr	6356	25430
x"00",	-- Hex Addr	6357	25431
x"00",	-- Hex Addr	6358	25432
x"00",	-- Hex Addr	6359	25433
x"00",	-- Hex Addr	635A	25434
x"00",	-- Hex Addr	635B	25435
x"00",	-- Hex Addr	635C	25436
x"00",	-- Hex Addr	635D	25437
x"00",	-- Hex Addr	635E	25438
x"00",	-- Hex Addr	635F	25439
x"00",	-- Hex Addr	6360	25440
x"00",	-- Hex Addr	6361	25441
x"00",	-- Hex Addr	6362	25442
x"00",	-- Hex Addr	6363	25443
x"00",	-- Hex Addr	6364	25444
x"00",	-- Hex Addr	6365	25445
x"00",	-- Hex Addr	6366	25446
x"00",	-- Hex Addr	6367	25447
x"00",	-- Hex Addr	6368	25448
x"00",	-- Hex Addr	6369	25449
x"00",	-- Hex Addr	636A	25450
x"00",	-- Hex Addr	636B	25451
x"00",	-- Hex Addr	636C	25452
x"00",	-- Hex Addr	636D	25453
x"00",	-- Hex Addr	636E	25454
x"00",	-- Hex Addr	636F	25455
x"00",	-- Hex Addr	6370	25456
x"00",	-- Hex Addr	6371	25457
x"00",	-- Hex Addr	6372	25458
x"00",	-- Hex Addr	6373	25459
x"00",	-- Hex Addr	6374	25460
x"00",	-- Hex Addr	6375	25461
x"00",	-- Hex Addr	6376	25462
x"00",	-- Hex Addr	6377	25463
x"00",	-- Hex Addr	6378	25464
x"00",	-- Hex Addr	6379	25465
x"00",	-- Hex Addr	637A	25466
x"00",	-- Hex Addr	637B	25467
x"00",	-- Hex Addr	637C	25468
x"00",	-- Hex Addr	637D	25469
x"00",	-- Hex Addr	637E	25470
x"00",	-- Hex Addr	637F	25471
x"00",	-- Hex Addr	6380	25472
x"00",	-- Hex Addr	6381	25473
x"00",	-- Hex Addr	6382	25474
x"00",	-- Hex Addr	6383	25475
x"00",	-- Hex Addr	6384	25476
x"00",	-- Hex Addr	6385	25477
x"00",	-- Hex Addr	6386	25478
x"00",	-- Hex Addr	6387	25479
x"00",	-- Hex Addr	6388	25480
x"00",	-- Hex Addr	6389	25481
x"00",	-- Hex Addr	638A	25482
x"00",	-- Hex Addr	638B	25483
x"00",	-- Hex Addr	638C	25484
x"00",	-- Hex Addr	638D	25485
x"00",	-- Hex Addr	638E	25486
x"00",	-- Hex Addr	638F	25487
x"00",	-- Hex Addr	6390	25488
x"00",	-- Hex Addr	6391	25489
x"00",	-- Hex Addr	6392	25490
x"00",	-- Hex Addr	6393	25491
x"00",	-- Hex Addr	6394	25492
x"00",	-- Hex Addr	6395	25493
x"00",	-- Hex Addr	6396	25494
x"00",	-- Hex Addr	6397	25495
x"00",	-- Hex Addr	6398	25496
x"00",	-- Hex Addr	6399	25497
x"00",	-- Hex Addr	639A	25498
x"00",	-- Hex Addr	639B	25499
x"00",	-- Hex Addr	639C	25500
x"00",	-- Hex Addr	639D	25501
x"00",	-- Hex Addr	639E	25502
x"00",	-- Hex Addr	639F	25503
x"00",	-- Hex Addr	63A0	25504
x"00",	-- Hex Addr	63A1	25505
x"00",	-- Hex Addr	63A2	25506
x"00",	-- Hex Addr	63A3	25507
x"00",	-- Hex Addr	63A4	25508
x"00",	-- Hex Addr	63A5	25509
x"00",	-- Hex Addr	63A6	25510
x"00",	-- Hex Addr	63A7	25511
x"00",	-- Hex Addr	63A8	25512
x"00",	-- Hex Addr	63A9	25513
x"00",	-- Hex Addr	63AA	25514
x"00",	-- Hex Addr	63AB	25515
x"00",	-- Hex Addr	63AC	25516
x"00",	-- Hex Addr	63AD	25517
x"00",	-- Hex Addr	63AE	25518
x"00",	-- Hex Addr	63AF	25519
x"00",	-- Hex Addr	63B0	25520
x"00",	-- Hex Addr	63B1	25521
x"00",	-- Hex Addr	63B2	25522
x"00",	-- Hex Addr	63B3	25523
x"00",	-- Hex Addr	63B4	25524
x"00",	-- Hex Addr	63B5	25525
x"00",	-- Hex Addr	63B6	25526
x"00",	-- Hex Addr	63B7	25527
x"00",	-- Hex Addr	63B8	25528
x"00",	-- Hex Addr	63B9	25529
x"00",	-- Hex Addr	63BA	25530
x"00",	-- Hex Addr	63BB	25531
x"00",	-- Hex Addr	63BC	25532
x"00",	-- Hex Addr	63BD	25533
x"00",	-- Hex Addr	63BE	25534
x"00",	-- Hex Addr	63BF	25535
x"00",	-- Hex Addr	63C0	25536
x"00",	-- Hex Addr	63C1	25537
x"00",	-- Hex Addr	63C2	25538
x"00",	-- Hex Addr	63C3	25539
x"00",	-- Hex Addr	63C4	25540
x"00",	-- Hex Addr	63C5	25541
x"00",	-- Hex Addr	63C6	25542
x"00",	-- Hex Addr	63C7	25543
x"00",	-- Hex Addr	63C8	25544
x"00",	-- Hex Addr	63C9	25545
x"00",	-- Hex Addr	63CA	25546
x"00",	-- Hex Addr	63CB	25547
x"00",	-- Hex Addr	63CC	25548
x"00",	-- Hex Addr	63CD	25549
x"00",	-- Hex Addr	63CE	25550
x"00",	-- Hex Addr	63CF	25551
x"00",	-- Hex Addr	63D0	25552
x"00",	-- Hex Addr	63D1	25553
x"00",	-- Hex Addr	63D2	25554
x"00",	-- Hex Addr	63D3	25555
x"00",	-- Hex Addr	63D4	25556
x"00",	-- Hex Addr	63D5	25557
x"00",	-- Hex Addr	63D6	25558
x"00",	-- Hex Addr	63D7	25559
x"00",	-- Hex Addr	63D8	25560
x"00",	-- Hex Addr	63D9	25561
x"00",	-- Hex Addr	63DA	25562
x"00",	-- Hex Addr	63DB	25563
x"00",	-- Hex Addr	63DC	25564
x"00",	-- Hex Addr	63DD	25565
x"00",	-- Hex Addr	63DE	25566
x"00",	-- Hex Addr	63DF	25567
x"00",	-- Hex Addr	63E0	25568
x"00",	-- Hex Addr	63E1	25569
x"00",	-- Hex Addr	63E2	25570
x"00",	-- Hex Addr	63E3	25571
x"00",	-- Hex Addr	63E4	25572
x"00",	-- Hex Addr	63E5	25573
x"00",	-- Hex Addr	63E6	25574
x"00",	-- Hex Addr	63E7	25575
x"00",	-- Hex Addr	63E8	25576
x"00",	-- Hex Addr	63E9	25577
x"00",	-- Hex Addr	63EA	25578
x"00",	-- Hex Addr	63EB	25579
x"00",	-- Hex Addr	63EC	25580
x"00",	-- Hex Addr	63ED	25581
x"00",	-- Hex Addr	63EE	25582
x"00",	-- Hex Addr	63EF	25583
x"00",	-- Hex Addr	63F0	25584
x"00",	-- Hex Addr	63F1	25585
x"00",	-- Hex Addr	63F2	25586
x"00",	-- Hex Addr	63F3	25587
x"00",	-- Hex Addr	63F4	25588
x"00",	-- Hex Addr	63F5	25589
x"00",	-- Hex Addr	63F6	25590
x"00",	-- Hex Addr	63F7	25591
x"00",	-- Hex Addr	63F8	25592
x"00",	-- Hex Addr	63F9	25593
x"00",	-- Hex Addr	63FA	25594
x"00",	-- Hex Addr	63FB	25595
x"00",	-- Hex Addr	63FC	25596
x"00",	-- Hex Addr	63FD	25597
x"00",	-- Hex Addr	63FE	25598
x"00",	-- Hex Addr	63FF	25599
x"00",	-- Hex Addr	6400	25600
x"00",	-- Hex Addr	6401	25601
x"00",	-- Hex Addr	6402	25602
x"00",	-- Hex Addr	6403	25603
x"00",	-- Hex Addr	6404	25604
x"00",	-- Hex Addr	6405	25605
x"00",	-- Hex Addr	6406	25606
x"00",	-- Hex Addr	6407	25607
x"00",	-- Hex Addr	6408	25608
x"00",	-- Hex Addr	6409	25609
x"00",	-- Hex Addr	640A	25610
x"00",	-- Hex Addr	640B	25611
x"00",	-- Hex Addr	640C	25612
x"00",	-- Hex Addr	640D	25613
x"00",	-- Hex Addr	640E	25614
x"00",	-- Hex Addr	640F	25615
x"00",	-- Hex Addr	6410	25616
x"00",	-- Hex Addr	6411	25617
x"00",	-- Hex Addr	6412	25618
x"00",	-- Hex Addr	6413	25619
x"00",	-- Hex Addr	6414	25620
x"00",	-- Hex Addr	6415	25621
x"00",	-- Hex Addr	6416	25622
x"00",	-- Hex Addr	6417	25623
x"00",	-- Hex Addr	6418	25624
x"00",	-- Hex Addr	6419	25625
x"00",	-- Hex Addr	641A	25626
x"00",	-- Hex Addr	641B	25627
x"00",	-- Hex Addr	641C	25628
x"00",	-- Hex Addr	641D	25629
x"00",	-- Hex Addr	641E	25630
x"00",	-- Hex Addr	641F	25631
x"00",	-- Hex Addr	6420	25632
x"00",	-- Hex Addr	6421	25633
x"00",	-- Hex Addr	6422	25634
x"00",	-- Hex Addr	6423	25635
x"00",	-- Hex Addr	6424	25636
x"00",	-- Hex Addr	6425	25637
x"00",	-- Hex Addr	6426	25638
x"00",	-- Hex Addr	6427	25639
x"00",	-- Hex Addr	6428	25640
x"00",	-- Hex Addr	6429	25641
x"00",	-- Hex Addr	642A	25642
x"00",	-- Hex Addr	642B	25643
x"00",	-- Hex Addr	642C	25644
x"00",	-- Hex Addr	642D	25645
x"00",	-- Hex Addr	642E	25646
x"00",	-- Hex Addr	642F	25647
x"00",	-- Hex Addr	6430	25648
x"00",	-- Hex Addr	6431	25649
x"00",	-- Hex Addr	6432	25650
x"00",	-- Hex Addr	6433	25651
x"00",	-- Hex Addr	6434	25652
x"00",	-- Hex Addr	6435	25653
x"00",	-- Hex Addr	6436	25654
x"00",	-- Hex Addr	6437	25655
x"00",	-- Hex Addr	6438	25656
x"00",	-- Hex Addr	6439	25657
x"00",	-- Hex Addr	643A	25658
x"00",	-- Hex Addr	643B	25659
x"00",	-- Hex Addr	643C	25660
x"00",	-- Hex Addr	643D	25661
x"00",	-- Hex Addr	643E	25662
x"00",	-- Hex Addr	643F	25663
x"00",	-- Hex Addr	6440	25664
x"00",	-- Hex Addr	6441	25665
x"00",	-- Hex Addr	6442	25666
x"00",	-- Hex Addr	6443	25667
x"00",	-- Hex Addr	6444	25668
x"00",	-- Hex Addr	6445	25669
x"00",	-- Hex Addr	6446	25670
x"00",	-- Hex Addr	6447	25671
x"00",	-- Hex Addr	6448	25672
x"00",	-- Hex Addr	6449	25673
x"00",	-- Hex Addr	644A	25674
x"00",	-- Hex Addr	644B	25675
x"00",	-- Hex Addr	644C	25676
x"00",	-- Hex Addr	644D	25677
x"00",	-- Hex Addr	644E	25678
x"00",	-- Hex Addr	644F	25679
x"00",	-- Hex Addr	6450	25680
x"00",	-- Hex Addr	6451	25681
x"00",	-- Hex Addr	6452	25682
x"00",	-- Hex Addr	6453	25683
x"00",	-- Hex Addr	6454	25684
x"00",	-- Hex Addr	6455	25685
x"00",	-- Hex Addr	6456	25686
x"00",	-- Hex Addr	6457	25687
x"00",	-- Hex Addr	6458	25688
x"00",	-- Hex Addr	6459	25689
x"00",	-- Hex Addr	645A	25690
x"00",	-- Hex Addr	645B	25691
x"00",	-- Hex Addr	645C	25692
x"00",	-- Hex Addr	645D	25693
x"00",	-- Hex Addr	645E	25694
x"00",	-- Hex Addr	645F	25695
x"00",	-- Hex Addr	6460	25696
x"00",	-- Hex Addr	6461	25697
x"00",	-- Hex Addr	6462	25698
x"00",	-- Hex Addr	6463	25699
x"00",	-- Hex Addr	6464	25700
x"00",	-- Hex Addr	6465	25701
x"00",	-- Hex Addr	6466	25702
x"00",	-- Hex Addr	6467	25703
x"00",	-- Hex Addr	6468	25704
x"00",	-- Hex Addr	6469	25705
x"00",	-- Hex Addr	646A	25706
x"00",	-- Hex Addr	646B	25707
x"00",	-- Hex Addr	646C	25708
x"00",	-- Hex Addr	646D	25709
x"00",	-- Hex Addr	646E	25710
x"00",	-- Hex Addr	646F	25711
x"00",	-- Hex Addr	6470	25712
x"00",	-- Hex Addr	6471	25713
x"00",	-- Hex Addr	6472	25714
x"00",	-- Hex Addr	6473	25715
x"00",	-- Hex Addr	6474	25716
x"00",	-- Hex Addr	6475	25717
x"00",	-- Hex Addr	6476	25718
x"00",	-- Hex Addr	6477	25719
x"00",	-- Hex Addr	6478	25720
x"00",	-- Hex Addr	6479	25721
x"00",	-- Hex Addr	647A	25722
x"00",	-- Hex Addr	647B	25723
x"00",	-- Hex Addr	647C	25724
x"00",	-- Hex Addr	647D	25725
x"00",	-- Hex Addr	647E	25726
x"00",	-- Hex Addr	647F	25727
x"00",	-- Hex Addr	6480	25728
x"00",	-- Hex Addr	6481	25729
x"00",	-- Hex Addr	6482	25730
x"00",	-- Hex Addr	6483	25731
x"00",	-- Hex Addr	6484	25732
x"00",	-- Hex Addr	6485	25733
x"00",	-- Hex Addr	6486	25734
x"00",	-- Hex Addr	6487	25735
x"00",	-- Hex Addr	6488	25736
x"00",	-- Hex Addr	6489	25737
x"00",	-- Hex Addr	648A	25738
x"00",	-- Hex Addr	648B	25739
x"00",	-- Hex Addr	648C	25740
x"00",	-- Hex Addr	648D	25741
x"00",	-- Hex Addr	648E	25742
x"00",	-- Hex Addr	648F	25743
x"00",	-- Hex Addr	6490	25744
x"00",	-- Hex Addr	6491	25745
x"00",	-- Hex Addr	6492	25746
x"00",	-- Hex Addr	6493	25747
x"00",	-- Hex Addr	6494	25748
x"00",	-- Hex Addr	6495	25749
x"00",	-- Hex Addr	6496	25750
x"00",	-- Hex Addr	6497	25751
x"00",	-- Hex Addr	6498	25752
x"00",	-- Hex Addr	6499	25753
x"00",	-- Hex Addr	649A	25754
x"00",	-- Hex Addr	649B	25755
x"00",	-- Hex Addr	649C	25756
x"00",	-- Hex Addr	649D	25757
x"00",	-- Hex Addr	649E	25758
x"00",	-- Hex Addr	649F	25759
x"00",	-- Hex Addr	64A0	25760
x"00",	-- Hex Addr	64A1	25761
x"00",	-- Hex Addr	64A2	25762
x"00",	-- Hex Addr	64A3	25763
x"00",	-- Hex Addr	64A4	25764
x"00",	-- Hex Addr	64A5	25765
x"00",	-- Hex Addr	64A6	25766
x"00",	-- Hex Addr	64A7	25767
x"00",	-- Hex Addr	64A8	25768
x"00",	-- Hex Addr	64A9	25769
x"00",	-- Hex Addr	64AA	25770
x"00",	-- Hex Addr	64AB	25771
x"00",	-- Hex Addr	64AC	25772
x"00",	-- Hex Addr	64AD	25773
x"00",	-- Hex Addr	64AE	25774
x"00",	-- Hex Addr	64AF	25775
x"00",	-- Hex Addr	64B0	25776
x"00",	-- Hex Addr	64B1	25777
x"00",	-- Hex Addr	64B2	25778
x"00",	-- Hex Addr	64B3	25779
x"00",	-- Hex Addr	64B4	25780
x"00",	-- Hex Addr	64B5	25781
x"00",	-- Hex Addr	64B6	25782
x"00",	-- Hex Addr	64B7	25783
x"00",	-- Hex Addr	64B8	25784
x"00",	-- Hex Addr	64B9	25785
x"00",	-- Hex Addr	64BA	25786
x"00",	-- Hex Addr	64BB	25787
x"00",	-- Hex Addr	64BC	25788
x"00",	-- Hex Addr	64BD	25789
x"00",	-- Hex Addr	64BE	25790
x"00",	-- Hex Addr	64BF	25791
x"00",	-- Hex Addr	64C0	25792
x"00",	-- Hex Addr	64C1	25793
x"00",	-- Hex Addr	64C2	25794
x"00",	-- Hex Addr	64C3	25795
x"00",	-- Hex Addr	64C4	25796
x"00",	-- Hex Addr	64C5	25797
x"00",	-- Hex Addr	64C6	25798
x"00",	-- Hex Addr	64C7	25799
x"00",	-- Hex Addr	64C8	25800
x"00",	-- Hex Addr	64C9	25801
x"00",	-- Hex Addr	64CA	25802
x"00",	-- Hex Addr	64CB	25803
x"00",	-- Hex Addr	64CC	25804
x"00",	-- Hex Addr	64CD	25805
x"00",	-- Hex Addr	64CE	25806
x"00",	-- Hex Addr	64CF	25807
x"00",	-- Hex Addr	64D0	25808
x"00",	-- Hex Addr	64D1	25809
x"00",	-- Hex Addr	64D2	25810
x"00",	-- Hex Addr	64D3	25811
x"00",	-- Hex Addr	64D4	25812
x"00",	-- Hex Addr	64D5	25813
x"00",	-- Hex Addr	64D6	25814
x"00",	-- Hex Addr	64D7	25815
x"00",	-- Hex Addr	64D8	25816
x"00",	-- Hex Addr	64D9	25817
x"00",	-- Hex Addr	64DA	25818
x"00",	-- Hex Addr	64DB	25819
x"00",	-- Hex Addr	64DC	25820
x"00",	-- Hex Addr	64DD	25821
x"00",	-- Hex Addr	64DE	25822
x"00",	-- Hex Addr	64DF	25823
x"00",	-- Hex Addr	64E0	25824
x"00",	-- Hex Addr	64E1	25825
x"00",	-- Hex Addr	64E2	25826
x"00",	-- Hex Addr	64E3	25827
x"00",	-- Hex Addr	64E4	25828
x"00",	-- Hex Addr	64E5	25829
x"00",	-- Hex Addr	64E6	25830
x"00",	-- Hex Addr	64E7	25831
x"00",	-- Hex Addr	64E8	25832
x"00",	-- Hex Addr	64E9	25833
x"00",	-- Hex Addr	64EA	25834
x"00",	-- Hex Addr	64EB	25835
x"00",	-- Hex Addr	64EC	25836
x"00",	-- Hex Addr	64ED	25837
x"00",	-- Hex Addr	64EE	25838
x"00",	-- Hex Addr	64EF	25839
x"00",	-- Hex Addr	64F0	25840
x"00",	-- Hex Addr	64F1	25841
x"00",	-- Hex Addr	64F2	25842
x"00",	-- Hex Addr	64F3	25843
x"00",	-- Hex Addr	64F4	25844
x"00",	-- Hex Addr	64F5	25845
x"00",	-- Hex Addr	64F6	25846
x"00",	-- Hex Addr	64F7	25847
x"00",	-- Hex Addr	64F8	25848
x"00",	-- Hex Addr	64F9	25849
x"00",	-- Hex Addr	64FA	25850
x"00",	-- Hex Addr	64FB	25851
x"00",	-- Hex Addr	64FC	25852
x"00",	-- Hex Addr	64FD	25853
x"00",	-- Hex Addr	64FE	25854
x"00",	-- Hex Addr	64FF	25855
x"00",	-- Hex Addr	6500	25856
x"00",	-- Hex Addr	6501	25857
x"00",	-- Hex Addr	6502	25858
x"00",	-- Hex Addr	6503	25859
x"00",	-- Hex Addr	6504	25860
x"00",	-- Hex Addr	6505	25861
x"00",	-- Hex Addr	6506	25862
x"00",	-- Hex Addr	6507	25863
x"00",	-- Hex Addr	6508	25864
x"00",	-- Hex Addr	6509	25865
x"00",	-- Hex Addr	650A	25866
x"00",	-- Hex Addr	650B	25867
x"00",	-- Hex Addr	650C	25868
x"00",	-- Hex Addr	650D	25869
x"00",	-- Hex Addr	650E	25870
x"00",	-- Hex Addr	650F	25871
x"00",	-- Hex Addr	6510	25872
x"00",	-- Hex Addr	6511	25873
x"00",	-- Hex Addr	6512	25874
x"00",	-- Hex Addr	6513	25875
x"00",	-- Hex Addr	6514	25876
x"00",	-- Hex Addr	6515	25877
x"00",	-- Hex Addr	6516	25878
x"00",	-- Hex Addr	6517	25879
x"00",	-- Hex Addr	6518	25880
x"00",	-- Hex Addr	6519	25881
x"00",	-- Hex Addr	651A	25882
x"00",	-- Hex Addr	651B	25883
x"00",	-- Hex Addr	651C	25884
x"00",	-- Hex Addr	651D	25885
x"00",	-- Hex Addr	651E	25886
x"00",	-- Hex Addr	651F	25887
x"00",	-- Hex Addr	6520	25888
x"00",	-- Hex Addr	6521	25889
x"00",	-- Hex Addr	6522	25890
x"00",	-- Hex Addr	6523	25891
x"00",	-- Hex Addr	6524	25892
x"00",	-- Hex Addr	6525	25893
x"00",	-- Hex Addr	6526	25894
x"00",	-- Hex Addr	6527	25895
x"00",	-- Hex Addr	6528	25896
x"00",	-- Hex Addr	6529	25897
x"00",	-- Hex Addr	652A	25898
x"00",	-- Hex Addr	652B	25899
x"00",	-- Hex Addr	652C	25900
x"00",	-- Hex Addr	652D	25901
x"00",	-- Hex Addr	652E	25902
x"00",	-- Hex Addr	652F	25903
x"00",	-- Hex Addr	6530	25904
x"00",	-- Hex Addr	6531	25905
x"00",	-- Hex Addr	6532	25906
x"00",	-- Hex Addr	6533	25907
x"00",	-- Hex Addr	6534	25908
x"00",	-- Hex Addr	6535	25909
x"00",	-- Hex Addr	6536	25910
x"00",	-- Hex Addr	6537	25911
x"00",	-- Hex Addr	6538	25912
x"00",	-- Hex Addr	6539	25913
x"00",	-- Hex Addr	653A	25914
x"00",	-- Hex Addr	653B	25915
x"00",	-- Hex Addr	653C	25916
x"00",	-- Hex Addr	653D	25917
x"00",	-- Hex Addr	653E	25918
x"00",	-- Hex Addr	653F	25919
x"00",	-- Hex Addr	6540	25920
x"00",	-- Hex Addr	6541	25921
x"00",	-- Hex Addr	6542	25922
x"00",	-- Hex Addr	6543	25923
x"00",	-- Hex Addr	6544	25924
x"00",	-- Hex Addr	6545	25925
x"00",	-- Hex Addr	6546	25926
x"00",	-- Hex Addr	6547	25927
x"00",	-- Hex Addr	6548	25928
x"00",	-- Hex Addr	6549	25929
x"00",	-- Hex Addr	654A	25930
x"00",	-- Hex Addr	654B	25931
x"00",	-- Hex Addr	654C	25932
x"00",	-- Hex Addr	654D	25933
x"00",	-- Hex Addr	654E	25934
x"00",	-- Hex Addr	654F	25935
x"00",	-- Hex Addr	6550	25936
x"00",	-- Hex Addr	6551	25937
x"00",	-- Hex Addr	6552	25938
x"00",	-- Hex Addr	6553	25939
x"00",	-- Hex Addr	6554	25940
x"00",	-- Hex Addr	6555	25941
x"00",	-- Hex Addr	6556	25942
x"00",	-- Hex Addr	6557	25943
x"00",	-- Hex Addr	6558	25944
x"00",	-- Hex Addr	6559	25945
x"00",	-- Hex Addr	655A	25946
x"00",	-- Hex Addr	655B	25947
x"00",	-- Hex Addr	655C	25948
x"00",	-- Hex Addr	655D	25949
x"00",	-- Hex Addr	655E	25950
x"00",	-- Hex Addr	655F	25951
x"00",	-- Hex Addr	6560	25952
x"00",	-- Hex Addr	6561	25953
x"00",	-- Hex Addr	6562	25954
x"00",	-- Hex Addr	6563	25955
x"00",	-- Hex Addr	6564	25956
x"00",	-- Hex Addr	6565	25957
x"00",	-- Hex Addr	6566	25958
x"00",	-- Hex Addr	6567	25959
x"00",	-- Hex Addr	6568	25960
x"00",	-- Hex Addr	6569	25961
x"00",	-- Hex Addr	656A	25962
x"00",	-- Hex Addr	656B	25963
x"00",	-- Hex Addr	656C	25964
x"00",	-- Hex Addr	656D	25965
x"00",	-- Hex Addr	656E	25966
x"00",	-- Hex Addr	656F	25967
x"00",	-- Hex Addr	6570	25968
x"00",	-- Hex Addr	6571	25969
x"00",	-- Hex Addr	6572	25970
x"00",	-- Hex Addr	6573	25971
x"00",	-- Hex Addr	6574	25972
x"00",	-- Hex Addr	6575	25973
x"00",	-- Hex Addr	6576	25974
x"00",	-- Hex Addr	6577	25975
x"00",	-- Hex Addr	6578	25976
x"00",	-- Hex Addr	6579	25977
x"00",	-- Hex Addr	657A	25978
x"00",	-- Hex Addr	657B	25979
x"00",	-- Hex Addr	657C	25980
x"00",	-- Hex Addr	657D	25981
x"00",	-- Hex Addr	657E	25982
x"00",	-- Hex Addr	657F	25983
x"00",	-- Hex Addr	6580	25984
x"00",	-- Hex Addr	6581	25985
x"00",	-- Hex Addr	6582	25986
x"00",	-- Hex Addr	6583	25987
x"00",	-- Hex Addr	6584	25988
x"00",	-- Hex Addr	6585	25989
x"00",	-- Hex Addr	6586	25990
x"00",	-- Hex Addr	6587	25991
x"00",	-- Hex Addr	6588	25992
x"00",	-- Hex Addr	6589	25993
x"00",	-- Hex Addr	658A	25994
x"00",	-- Hex Addr	658B	25995
x"00",	-- Hex Addr	658C	25996
x"00",	-- Hex Addr	658D	25997
x"00",	-- Hex Addr	658E	25998
x"00",	-- Hex Addr	658F	25999
x"00",	-- Hex Addr	6590	26000
x"00",	-- Hex Addr	6591	26001
x"00",	-- Hex Addr	6592	26002
x"00",	-- Hex Addr	6593	26003
x"00",	-- Hex Addr	6594	26004
x"00",	-- Hex Addr	6595	26005
x"00",	-- Hex Addr	6596	26006
x"00",	-- Hex Addr	6597	26007
x"00",	-- Hex Addr	6598	26008
x"00",	-- Hex Addr	6599	26009
x"00",	-- Hex Addr	659A	26010
x"00",	-- Hex Addr	659B	26011
x"00",	-- Hex Addr	659C	26012
x"00",	-- Hex Addr	659D	26013
x"00",	-- Hex Addr	659E	26014
x"00",	-- Hex Addr	659F	26015
x"00",	-- Hex Addr	65A0	26016
x"00",	-- Hex Addr	65A1	26017
x"00",	-- Hex Addr	65A2	26018
x"00",	-- Hex Addr	65A3	26019
x"00",	-- Hex Addr	65A4	26020
x"00",	-- Hex Addr	65A5	26021
x"00",	-- Hex Addr	65A6	26022
x"00",	-- Hex Addr	65A7	26023
x"00",	-- Hex Addr	65A8	26024
x"00",	-- Hex Addr	65A9	26025
x"00",	-- Hex Addr	65AA	26026
x"00",	-- Hex Addr	65AB	26027
x"00",	-- Hex Addr	65AC	26028
x"00",	-- Hex Addr	65AD	26029
x"00",	-- Hex Addr	65AE	26030
x"00",	-- Hex Addr	65AF	26031
x"00",	-- Hex Addr	65B0	26032
x"00",	-- Hex Addr	65B1	26033
x"00",	-- Hex Addr	65B2	26034
x"00",	-- Hex Addr	65B3	26035
x"00",	-- Hex Addr	65B4	26036
x"00",	-- Hex Addr	65B5	26037
x"00",	-- Hex Addr	65B6	26038
x"00",	-- Hex Addr	65B7	26039
x"00",	-- Hex Addr	65B8	26040
x"00",	-- Hex Addr	65B9	26041
x"00",	-- Hex Addr	65BA	26042
x"00",	-- Hex Addr	65BB	26043
x"00",	-- Hex Addr	65BC	26044
x"00",	-- Hex Addr	65BD	26045
x"00",	-- Hex Addr	65BE	26046
x"00",	-- Hex Addr	65BF	26047
x"00",	-- Hex Addr	65C0	26048
x"00",	-- Hex Addr	65C1	26049
x"00",	-- Hex Addr	65C2	26050
x"00",	-- Hex Addr	65C3	26051
x"00",	-- Hex Addr	65C4	26052
x"00",	-- Hex Addr	65C5	26053
x"00",	-- Hex Addr	65C6	26054
x"00",	-- Hex Addr	65C7	26055
x"00",	-- Hex Addr	65C8	26056
x"00",	-- Hex Addr	65C9	26057
x"00",	-- Hex Addr	65CA	26058
x"00",	-- Hex Addr	65CB	26059
x"00",	-- Hex Addr	65CC	26060
x"00",	-- Hex Addr	65CD	26061
x"00",	-- Hex Addr	65CE	26062
x"00",	-- Hex Addr	65CF	26063
x"00",	-- Hex Addr	65D0	26064
x"00",	-- Hex Addr	65D1	26065
x"00",	-- Hex Addr	65D2	26066
x"00",	-- Hex Addr	65D3	26067
x"00",	-- Hex Addr	65D4	26068
x"00",	-- Hex Addr	65D5	26069
x"00",	-- Hex Addr	65D6	26070
x"00",	-- Hex Addr	65D7	26071
x"00",	-- Hex Addr	65D8	26072
x"00",	-- Hex Addr	65D9	26073
x"00",	-- Hex Addr	65DA	26074
x"00",	-- Hex Addr	65DB	26075
x"00",	-- Hex Addr	65DC	26076
x"00",	-- Hex Addr	65DD	26077
x"00",	-- Hex Addr	65DE	26078
x"00",	-- Hex Addr	65DF	26079
x"00",	-- Hex Addr	65E0	26080
x"00",	-- Hex Addr	65E1	26081
x"00",	-- Hex Addr	65E2	26082
x"00",	-- Hex Addr	65E3	26083
x"00",	-- Hex Addr	65E4	26084
x"00",	-- Hex Addr	65E5	26085
x"00",	-- Hex Addr	65E6	26086
x"00",	-- Hex Addr	65E7	26087
x"00",	-- Hex Addr	65E8	26088
x"00",	-- Hex Addr	65E9	26089
x"00",	-- Hex Addr	65EA	26090
x"00",	-- Hex Addr	65EB	26091
x"00",	-- Hex Addr	65EC	26092
x"00",	-- Hex Addr	65ED	26093
x"00",	-- Hex Addr	65EE	26094
x"00",	-- Hex Addr	65EF	26095
x"00",	-- Hex Addr	65F0	26096
x"00",	-- Hex Addr	65F1	26097
x"00",	-- Hex Addr	65F2	26098
x"00",	-- Hex Addr	65F3	26099
x"00",	-- Hex Addr	65F4	26100
x"00",	-- Hex Addr	65F5	26101
x"00",	-- Hex Addr	65F6	26102
x"00",	-- Hex Addr	65F7	26103
x"00",	-- Hex Addr	65F8	26104
x"00",	-- Hex Addr	65F9	26105
x"00",	-- Hex Addr	65FA	26106
x"00",	-- Hex Addr	65FB	26107
x"00",	-- Hex Addr	65FC	26108
x"00",	-- Hex Addr	65FD	26109
x"00",	-- Hex Addr	65FE	26110
x"00",	-- Hex Addr	65FF	26111
x"00",	-- Hex Addr	6600	26112
x"00",	-- Hex Addr	6601	26113
x"00",	-- Hex Addr	6602	26114
x"00",	-- Hex Addr	6603	26115
x"00",	-- Hex Addr	6604	26116
x"00",	-- Hex Addr	6605	26117
x"00",	-- Hex Addr	6606	26118
x"00",	-- Hex Addr	6607	26119
x"00",	-- Hex Addr	6608	26120
x"00",	-- Hex Addr	6609	26121
x"00",	-- Hex Addr	660A	26122
x"00",	-- Hex Addr	660B	26123
x"00",	-- Hex Addr	660C	26124
x"00",	-- Hex Addr	660D	26125
x"00",	-- Hex Addr	660E	26126
x"00",	-- Hex Addr	660F	26127
x"00",	-- Hex Addr	6610	26128
x"00",	-- Hex Addr	6611	26129
x"00",	-- Hex Addr	6612	26130
x"00",	-- Hex Addr	6613	26131
x"00",	-- Hex Addr	6614	26132
x"00",	-- Hex Addr	6615	26133
x"00",	-- Hex Addr	6616	26134
x"00",	-- Hex Addr	6617	26135
x"00",	-- Hex Addr	6618	26136
x"00",	-- Hex Addr	6619	26137
x"00",	-- Hex Addr	661A	26138
x"00",	-- Hex Addr	661B	26139
x"00",	-- Hex Addr	661C	26140
x"00",	-- Hex Addr	661D	26141
x"00",	-- Hex Addr	661E	26142
x"00",	-- Hex Addr	661F	26143
x"00",	-- Hex Addr	6620	26144
x"00",	-- Hex Addr	6621	26145
x"00",	-- Hex Addr	6622	26146
x"00",	-- Hex Addr	6623	26147
x"00",	-- Hex Addr	6624	26148
x"00",	-- Hex Addr	6625	26149
x"00",	-- Hex Addr	6626	26150
x"00",	-- Hex Addr	6627	26151
x"00",	-- Hex Addr	6628	26152
x"00",	-- Hex Addr	6629	26153
x"00",	-- Hex Addr	662A	26154
x"00",	-- Hex Addr	662B	26155
x"00",	-- Hex Addr	662C	26156
x"00",	-- Hex Addr	662D	26157
x"00",	-- Hex Addr	662E	26158
x"00",	-- Hex Addr	662F	26159
x"00",	-- Hex Addr	6630	26160
x"00",	-- Hex Addr	6631	26161
x"00",	-- Hex Addr	6632	26162
x"00",	-- Hex Addr	6633	26163
x"00",	-- Hex Addr	6634	26164
x"00",	-- Hex Addr	6635	26165
x"00",	-- Hex Addr	6636	26166
x"00",	-- Hex Addr	6637	26167
x"00",	-- Hex Addr	6638	26168
x"00",	-- Hex Addr	6639	26169
x"00",	-- Hex Addr	663A	26170
x"00",	-- Hex Addr	663B	26171
x"00",	-- Hex Addr	663C	26172
x"00",	-- Hex Addr	663D	26173
x"00",	-- Hex Addr	663E	26174
x"00",	-- Hex Addr	663F	26175
x"00",	-- Hex Addr	6640	26176
x"00",	-- Hex Addr	6641	26177
x"00",	-- Hex Addr	6642	26178
x"00",	-- Hex Addr	6643	26179
x"00",	-- Hex Addr	6644	26180
x"00",	-- Hex Addr	6645	26181
x"00",	-- Hex Addr	6646	26182
x"00",	-- Hex Addr	6647	26183
x"00",	-- Hex Addr	6648	26184
x"00",	-- Hex Addr	6649	26185
x"00",	-- Hex Addr	664A	26186
x"00",	-- Hex Addr	664B	26187
x"00",	-- Hex Addr	664C	26188
x"00",	-- Hex Addr	664D	26189
x"00",	-- Hex Addr	664E	26190
x"00",	-- Hex Addr	664F	26191
x"00",	-- Hex Addr	6650	26192
x"00",	-- Hex Addr	6651	26193
x"00",	-- Hex Addr	6652	26194
x"00",	-- Hex Addr	6653	26195
x"00",	-- Hex Addr	6654	26196
x"00",	-- Hex Addr	6655	26197
x"00",	-- Hex Addr	6656	26198
x"00",	-- Hex Addr	6657	26199
x"00",	-- Hex Addr	6658	26200
x"00",	-- Hex Addr	6659	26201
x"00",	-- Hex Addr	665A	26202
x"00",	-- Hex Addr	665B	26203
x"00",	-- Hex Addr	665C	26204
x"00",	-- Hex Addr	665D	26205
x"00",	-- Hex Addr	665E	26206
x"00",	-- Hex Addr	665F	26207
x"00",	-- Hex Addr	6660	26208
x"00",	-- Hex Addr	6661	26209
x"00",	-- Hex Addr	6662	26210
x"00",	-- Hex Addr	6663	26211
x"00",	-- Hex Addr	6664	26212
x"00",	-- Hex Addr	6665	26213
x"00",	-- Hex Addr	6666	26214
x"00",	-- Hex Addr	6667	26215
x"00",	-- Hex Addr	6668	26216
x"00",	-- Hex Addr	6669	26217
x"00",	-- Hex Addr	666A	26218
x"00",	-- Hex Addr	666B	26219
x"00",	-- Hex Addr	666C	26220
x"00",	-- Hex Addr	666D	26221
x"00",	-- Hex Addr	666E	26222
x"00",	-- Hex Addr	666F	26223
x"00",	-- Hex Addr	6670	26224
x"00",	-- Hex Addr	6671	26225
x"00",	-- Hex Addr	6672	26226
x"00",	-- Hex Addr	6673	26227
x"00",	-- Hex Addr	6674	26228
x"00",	-- Hex Addr	6675	26229
x"00",	-- Hex Addr	6676	26230
x"00",	-- Hex Addr	6677	26231
x"00",	-- Hex Addr	6678	26232
x"00",	-- Hex Addr	6679	26233
x"00",	-- Hex Addr	667A	26234
x"00",	-- Hex Addr	667B	26235
x"00",	-- Hex Addr	667C	26236
x"00",	-- Hex Addr	667D	26237
x"00",	-- Hex Addr	667E	26238
x"00",	-- Hex Addr	667F	26239
x"00",	-- Hex Addr	6680	26240
x"00",	-- Hex Addr	6681	26241
x"00",	-- Hex Addr	6682	26242
x"00",	-- Hex Addr	6683	26243
x"00",	-- Hex Addr	6684	26244
x"00",	-- Hex Addr	6685	26245
x"00",	-- Hex Addr	6686	26246
x"00",	-- Hex Addr	6687	26247
x"00",	-- Hex Addr	6688	26248
x"00",	-- Hex Addr	6689	26249
x"00",	-- Hex Addr	668A	26250
x"00",	-- Hex Addr	668B	26251
x"00",	-- Hex Addr	668C	26252
x"00",	-- Hex Addr	668D	26253
x"00",	-- Hex Addr	668E	26254
x"00",	-- Hex Addr	668F	26255
x"00",	-- Hex Addr	6690	26256
x"00",	-- Hex Addr	6691	26257
x"00",	-- Hex Addr	6692	26258
x"00",	-- Hex Addr	6693	26259
x"00",	-- Hex Addr	6694	26260
x"00",	-- Hex Addr	6695	26261
x"00",	-- Hex Addr	6696	26262
x"00",	-- Hex Addr	6697	26263
x"00",	-- Hex Addr	6698	26264
x"00",	-- Hex Addr	6699	26265
x"00",	-- Hex Addr	669A	26266
x"00",	-- Hex Addr	669B	26267
x"00",	-- Hex Addr	669C	26268
x"00",	-- Hex Addr	669D	26269
x"00",	-- Hex Addr	669E	26270
x"00",	-- Hex Addr	669F	26271
x"00",	-- Hex Addr	66A0	26272
x"00",	-- Hex Addr	66A1	26273
x"00",	-- Hex Addr	66A2	26274
x"00",	-- Hex Addr	66A3	26275
x"00",	-- Hex Addr	66A4	26276
x"00",	-- Hex Addr	66A5	26277
x"00",	-- Hex Addr	66A6	26278
x"00",	-- Hex Addr	66A7	26279
x"00",	-- Hex Addr	66A8	26280
x"00",	-- Hex Addr	66A9	26281
x"00",	-- Hex Addr	66AA	26282
x"00",	-- Hex Addr	66AB	26283
x"00",	-- Hex Addr	66AC	26284
x"00",	-- Hex Addr	66AD	26285
x"00",	-- Hex Addr	66AE	26286
x"00",	-- Hex Addr	66AF	26287
x"00",	-- Hex Addr	66B0	26288
x"00",	-- Hex Addr	66B1	26289
x"00",	-- Hex Addr	66B2	26290
x"00",	-- Hex Addr	66B3	26291
x"00",	-- Hex Addr	66B4	26292
x"00",	-- Hex Addr	66B5	26293
x"00",	-- Hex Addr	66B6	26294
x"00",	-- Hex Addr	66B7	26295
x"00",	-- Hex Addr	66B8	26296
x"00",	-- Hex Addr	66B9	26297
x"00",	-- Hex Addr	66BA	26298
x"00",	-- Hex Addr	66BB	26299
x"00",	-- Hex Addr	66BC	26300
x"00",	-- Hex Addr	66BD	26301
x"00",	-- Hex Addr	66BE	26302
x"00",	-- Hex Addr	66BF	26303
x"00",	-- Hex Addr	66C0	26304
x"00",	-- Hex Addr	66C1	26305
x"00",	-- Hex Addr	66C2	26306
x"00",	-- Hex Addr	66C3	26307
x"00",	-- Hex Addr	66C4	26308
x"00",	-- Hex Addr	66C5	26309
x"00",	-- Hex Addr	66C6	26310
x"00",	-- Hex Addr	66C7	26311
x"00",	-- Hex Addr	66C8	26312
x"00",	-- Hex Addr	66C9	26313
x"00",	-- Hex Addr	66CA	26314
x"00",	-- Hex Addr	66CB	26315
x"00",	-- Hex Addr	66CC	26316
x"00",	-- Hex Addr	66CD	26317
x"00",	-- Hex Addr	66CE	26318
x"00",	-- Hex Addr	66CF	26319
x"00",	-- Hex Addr	66D0	26320
x"00",	-- Hex Addr	66D1	26321
x"00",	-- Hex Addr	66D2	26322
x"00",	-- Hex Addr	66D3	26323
x"00",	-- Hex Addr	66D4	26324
x"00",	-- Hex Addr	66D5	26325
x"00",	-- Hex Addr	66D6	26326
x"00",	-- Hex Addr	66D7	26327
x"00",	-- Hex Addr	66D8	26328
x"00",	-- Hex Addr	66D9	26329
x"00",	-- Hex Addr	66DA	26330
x"00",	-- Hex Addr	66DB	26331
x"00",	-- Hex Addr	66DC	26332
x"00",	-- Hex Addr	66DD	26333
x"00",	-- Hex Addr	66DE	26334
x"00",	-- Hex Addr	66DF	26335
x"00",	-- Hex Addr	66E0	26336
x"00",	-- Hex Addr	66E1	26337
x"00",	-- Hex Addr	66E2	26338
x"00",	-- Hex Addr	66E3	26339
x"00",	-- Hex Addr	66E4	26340
x"00",	-- Hex Addr	66E5	26341
x"00",	-- Hex Addr	66E6	26342
x"00",	-- Hex Addr	66E7	26343
x"00",	-- Hex Addr	66E8	26344
x"00",	-- Hex Addr	66E9	26345
x"00",	-- Hex Addr	66EA	26346
x"00",	-- Hex Addr	66EB	26347
x"00",	-- Hex Addr	66EC	26348
x"00",	-- Hex Addr	66ED	26349
x"00",	-- Hex Addr	66EE	26350
x"00",	-- Hex Addr	66EF	26351
x"00",	-- Hex Addr	66F0	26352
x"00",	-- Hex Addr	66F1	26353
x"00",	-- Hex Addr	66F2	26354
x"00",	-- Hex Addr	66F3	26355
x"00",	-- Hex Addr	66F4	26356
x"00",	-- Hex Addr	66F5	26357
x"00",	-- Hex Addr	66F6	26358
x"00",	-- Hex Addr	66F7	26359
x"00",	-- Hex Addr	66F8	26360
x"00",	-- Hex Addr	66F9	26361
x"00",	-- Hex Addr	66FA	26362
x"00",	-- Hex Addr	66FB	26363
x"00",	-- Hex Addr	66FC	26364
x"00",	-- Hex Addr	66FD	26365
x"00",	-- Hex Addr	66FE	26366
x"00",	-- Hex Addr	66FF	26367
x"00",	-- Hex Addr	6700	26368
x"00",	-- Hex Addr	6701	26369
x"00",	-- Hex Addr	6702	26370
x"00",	-- Hex Addr	6703	26371
x"00",	-- Hex Addr	6704	26372
x"00",	-- Hex Addr	6705	26373
x"00",	-- Hex Addr	6706	26374
x"00",	-- Hex Addr	6707	26375
x"00",	-- Hex Addr	6708	26376
x"00",	-- Hex Addr	6709	26377
x"00",	-- Hex Addr	670A	26378
x"00",	-- Hex Addr	670B	26379
x"00",	-- Hex Addr	670C	26380
x"00",	-- Hex Addr	670D	26381
x"00",	-- Hex Addr	670E	26382
x"00",	-- Hex Addr	670F	26383
x"00",	-- Hex Addr	6710	26384
x"00",	-- Hex Addr	6711	26385
x"00",	-- Hex Addr	6712	26386
x"00",	-- Hex Addr	6713	26387
x"00",	-- Hex Addr	6714	26388
x"00",	-- Hex Addr	6715	26389
x"00",	-- Hex Addr	6716	26390
x"00",	-- Hex Addr	6717	26391
x"00",	-- Hex Addr	6718	26392
x"00",	-- Hex Addr	6719	26393
x"00",	-- Hex Addr	671A	26394
x"00",	-- Hex Addr	671B	26395
x"00",	-- Hex Addr	671C	26396
x"00",	-- Hex Addr	671D	26397
x"00",	-- Hex Addr	671E	26398
x"00",	-- Hex Addr	671F	26399
x"00",	-- Hex Addr	6720	26400
x"00",	-- Hex Addr	6721	26401
x"00",	-- Hex Addr	6722	26402
x"00",	-- Hex Addr	6723	26403
x"00",	-- Hex Addr	6724	26404
x"00",	-- Hex Addr	6725	26405
x"00",	-- Hex Addr	6726	26406
x"00",	-- Hex Addr	6727	26407
x"00",	-- Hex Addr	6728	26408
x"00",	-- Hex Addr	6729	26409
x"00",	-- Hex Addr	672A	26410
x"00",	-- Hex Addr	672B	26411
x"00",	-- Hex Addr	672C	26412
x"00",	-- Hex Addr	672D	26413
x"00",	-- Hex Addr	672E	26414
x"00",	-- Hex Addr	672F	26415
x"00",	-- Hex Addr	6730	26416
x"00",	-- Hex Addr	6731	26417
x"00",	-- Hex Addr	6732	26418
x"00",	-- Hex Addr	6733	26419
x"00",	-- Hex Addr	6734	26420
x"00",	-- Hex Addr	6735	26421
x"00",	-- Hex Addr	6736	26422
x"00",	-- Hex Addr	6737	26423
x"00",	-- Hex Addr	6738	26424
x"00",	-- Hex Addr	6739	26425
x"00",	-- Hex Addr	673A	26426
x"00",	-- Hex Addr	673B	26427
x"00",	-- Hex Addr	673C	26428
x"00",	-- Hex Addr	673D	26429
x"00",	-- Hex Addr	673E	26430
x"00",	-- Hex Addr	673F	26431
x"00",	-- Hex Addr	6740	26432
x"00",	-- Hex Addr	6741	26433
x"00",	-- Hex Addr	6742	26434
x"00",	-- Hex Addr	6743	26435
x"00",	-- Hex Addr	6744	26436
x"00",	-- Hex Addr	6745	26437
x"00",	-- Hex Addr	6746	26438
x"00",	-- Hex Addr	6747	26439
x"00",	-- Hex Addr	6748	26440
x"00",	-- Hex Addr	6749	26441
x"00",	-- Hex Addr	674A	26442
x"00",	-- Hex Addr	674B	26443
x"00",	-- Hex Addr	674C	26444
x"00",	-- Hex Addr	674D	26445
x"00",	-- Hex Addr	674E	26446
x"00",	-- Hex Addr	674F	26447
x"00",	-- Hex Addr	6750	26448
x"00",	-- Hex Addr	6751	26449
x"00",	-- Hex Addr	6752	26450
x"00",	-- Hex Addr	6753	26451
x"00",	-- Hex Addr	6754	26452
x"00",	-- Hex Addr	6755	26453
x"00",	-- Hex Addr	6756	26454
x"00",	-- Hex Addr	6757	26455
x"00",	-- Hex Addr	6758	26456
x"00",	-- Hex Addr	6759	26457
x"00",	-- Hex Addr	675A	26458
x"00",	-- Hex Addr	675B	26459
x"00",	-- Hex Addr	675C	26460
x"00",	-- Hex Addr	675D	26461
x"00",	-- Hex Addr	675E	26462
x"00",	-- Hex Addr	675F	26463
x"00",	-- Hex Addr	6760	26464
x"00",	-- Hex Addr	6761	26465
x"00",	-- Hex Addr	6762	26466
x"00",	-- Hex Addr	6763	26467
x"00",	-- Hex Addr	6764	26468
x"00",	-- Hex Addr	6765	26469
x"00",	-- Hex Addr	6766	26470
x"00",	-- Hex Addr	6767	26471
x"00",	-- Hex Addr	6768	26472
x"00",	-- Hex Addr	6769	26473
x"00",	-- Hex Addr	676A	26474
x"00",	-- Hex Addr	676B	26475
x"00",	-- Hex Addr	676C	26476
x"00",	-- Hex Addr	676D	26477
x"00",	-- Hex Addr	676E	26478
x"00",	-- Hex Addr	676F	26479
x"00",	-- Hex Addr	6770	26480
x"00",	-- Hex Addr	6771	26481
x"00",	-- Hex Addr	6772	26482
x"00",	-- Hex Addr	6773	26483
x"00",	-- Hex Addr	6774	26484
x"00",	-- Hex Addr	6775	26485
x"00",	-- Hex Addr	6776	26486
x"00",	-- Hex Addr	6777	26487
x"00",	-- Hex Addr	6778	26488
x"00",	-- Hex Addr	6779	26489
x"00",	-- Hex Addr	677A	26490
x"00",	-- Hex Addr	677B	26491
x"00",	-- Hex Addr	677C	26492
x"00",	-- Hex Addr	677D	26493
x"00",	-- Hex Addr	677E	26494
x"00",	-- Hex Addr	677F	26495
x"00",	-- Hex Addr	6780	26496
x"00",	-- Hex Addr	6781	26497
x"00",	-- Hex Addr	6782	26498
x"00",	-- Hex Addr	6783	26499
x"00",	-- Hex Addr	6784	26500
x"00",	-- Hex Addr	6785	26501
x"00",	-- Hex Addr	6786	26502
x"00",	-- Hex Addr	6787	26503
x"00",	-- Hex Addr	6788	26504
x"00",	-- Hex Addr	6789	26505
x"00",	-- Hex Addr	678A	26506
x"00",	-- Hex Addr	678B	26507
x"00",	-- Hex Addr	678C	26508
x"00",	-- Hex Addr	678D	26509
x"00",	-- Hex Addr	678E	26510
x"00",	-- Hex Addr	678F	26511
x"00",	-- Hex Addr	6790	26512
x"00",	-- Hex Addr	6791	26513
x"00",	-- Hex Addr	6792	26514
x"00",	-- Hex Addr	6793	26515
x"00",	-- Hex Addr	6794	26516
x"00",	-- Hex Addr	6795	26517
x"00",	-- Hex Addr	6796	26518
x"00",	-- Hex Addr	6797	26519
x"00",	-- Hex Addr	6798	26520
x"00",	-- Hex Addr	6799	26521
x"00",	-- Hex Addr	679A	26522
x"00",	-- Hex Addr	679B	26523
x"00",	-- Hex Addr	679C	26524
x"00",	-- Hex Addr	679D	26525
x"00",	-- Hex Addr	679E	26526
x"00",	-- Hex Addr	679F	26527
x"00",	-- Hex Addr	67A0	26528
x"00",	-- Hex Addr	67A1	26529
x"00",	-- Hex Addr	67A2	26530
x"00",	-- Hex Addr	67A3	26531
x"00",	-- Hex Addr	67A4	26532
x"00",	-- Hex Addr	67A5	26533
x"00",	-- Hex Addr	67A6	26534
x"00",	-- Hex Addr	67A7	26535
x"00",	-- Hex Addr	67A8	26536
x"00",	-- Hex Addr	67A9	26537
x"00",	-- Hex Addr	67AA	26538
x"00",	-- Hex Addr	67AB	26539
x"00",	-- Hex Addr	67AC	26540
x"00",	-- Hex Addr	67AD	26541
x"00",	-- Hex Addr	67AE	26542
x"00",	-- Hex Addr	67AF	26543
x"00",	-- Hex Addr	67B0	26544
x"00",	-- Hex Addr	67B1	26545
x"00",	-- Hex Addr	67B2	26546
x"00",	-- Hex Addr	67B3	26547
x"00",	-- Hex Addr	67B4	26548
x"00",	-- Hex Addr	67B5	26549
x"00",	-- Hex Addr	67B6	26550
x"00",	-- Hex Addr	67B7	26551
x"00",	-- Hex Addr	67B8	26552
x"00",	-- Hex Addr	67B9	26553
x"00",	-- Hex Addr	67BA	26554
x"00",	-- Hex Addr	67BB	26555
x"00",	-- Hex Addr	67BC	26556
x"00",	-- Hex Addr	67BD	26557
x"00",	-- Hex Addr	67BE	26558
x"00",	-- Hex Addr	67BF	26559
x"00",	-- Hex Addr	67C0	26560
x"00",	-- Hex Addr	67C1	26561
x"00",	-- Hex Addr	67C2	26562
x"00",	-- Hex Addr	67C3	26563
x"00",	-- Hex Addr	67C4	26564
x"00",	-- Hex Addr	67C5	26565
x"00",	-- Hex Addr	67C6	26566
x"00",	-- Hex Addr	67C7	26567
x"00",	-- Hex Addr	67C8	26568
x"00",	-- Hex Addr	67C9	26569
x"00",	-- Hex Addr	67CA	26570
x"00",	-- Hex Addr	67CB	26571
x"00",	-- Hex Addr	67CC	26572
x"00",	-- Hex Addr	67CD	26573
x"00",	-- Hex Addr	67CE	26574
x"00",	-- Hex Addr	67CF	26575
x"00",	-- Hex Addr	67D0	26576
x"00",	-- Hex Addr	67D1	26577
x"00",	-- Hex Addr	67D2	26578
x"00",	-- Hex Addr	67D3	26579
x"00",	-- Hex Addr	67D4	26580
x"00",	-- Hex Addr	67D5	26581
x"00",	-- Hex Addr	67D6	26582
x"00",	-- Hex Addr	67D7	26583
x"00",	-- Hex Addr	67D8	26584
x"00",	-- Hex Addr	67D9	26585
x"00",	-- Hex Addr	67DA	26586
x"00",	-- Hex Addr	67DB	26587
x"00",	-- Hex Addr	67DC	26588
x"00",	-- Hex Addr	67DD	26589
x"00",	-- Hex Addr	67DE	26590
x"00",	-- Hex Addr	67DF	26591
x"00",	-- Hex Addr	67E0	26592
x"00",	-- Hex Addr	67E1	26593
x"00",	-- Hex Addr	67E2	26594
x"00",	-- Hex Addr	67E3	26595
x"00",	-- Hex Addr	67E4	26596
x"00",	-- Hex Addr	67E5	26597
x"00",	-- Hex Addr	67E6	26598
x"00",	-- Hex Addr	67E7	26599
x"00",	-- Hex Addr	67E8	26600
x"00",	-- Hex Addr	67E9	26601
x"00",	-- Hex Addr	67EA	26602
x"00",	-- Hex Addr	67EB	26603
x"00",	-- Hex Addr	67EC	26604
x"00",	-- Hex Addr	67ED	26605
x"00",	-- Hex Addr	67EE	26606
x"00",	-- Hex Addr	67EF	26607
x"00",	-- Hex Addr	67F0	26608
x"00",	-- Hex Addr	67F1	26609
x"00",	-- Hex Addr	67F2	26610
x"00",	-- Hex Addr	67F3	26611
x"00",	-- Hex Addr	67F4	26612
x"00",	-- Hex Addr	67F5	26613
x"00",	-- Hex Addr	67F6	26614
x"00",	-- Hex Addr	67F7	26615
x"00",	-- Hex Addr	67F8	26616
x"00",	-- Hex Addr	67F9	26617
x"00",	-- Hex Addr	67FA	26618
x"00",	-- Hex Addr	67FB	26619
x"00",	-- Hex Addr	67FC	26620
x"00",	-- Hex Addr	67FD	26621
x"00",	-- Hex Addr	67FE	26622
x"00",	-- Hex Addr	67FF	26623
x"00",	-- Hex Addr	6800	26624
x"00",	-- Hex Addr	6801	26625
x"00",	-- Hex Addr	6802	26626
x"00",	-- Hex Addr	6803	26627
x"00",	-- Hex Addr	6804	26628
x"00",	-- Hex Addr	6805	26629
x"00",	-- Hex Addr	6806	26630
x"00",	-- Hex Addr	6807	26631
x"00",	-- Hex Addr	6808	26632
x"00",	-- Hex Addr	6809	26633
x"00",	-- Hex Addr	680A	26634
x"00",	-- Hex Addr	680B	26635
x"00",	-- Hex Addr	680C	26636
x"00",	-- Hex Addr	680D	26637
x"00",	-- Hex Addr	680E	26638
x"00",	-- Hex Addr	680F	26639
x"00",	-- Hex Addr	6810	26640
x"00",	-- Hex Addr	6811	26641
x"00",	-- Hex Addr	6812	26642
x"00",	-- Hex Addr	6813	26643
x"00",	-- Hex Addr	6814	26644
x"00",	-- Hex Addr	6815	26645
x"00",	-- Hex Addr	6816	26646
x"00",	-- Hex Addr	6817	26647
x"00",	-- Hex Addr	6818	26648
x"00",	-- Hex Addr	6819	26649
x"00",	-- Hex Addr	681A	26650
x"00",	-- Hex Addr	681B	26651
x"00",	-- Hex Addr	681C	26652
x"00",	-- Hex Addr	681D	26653
x"00",	-- Hex Addr	681E	26654
x"00",	-- Hex Addr	681F	26655
x"00",	-- Hex Addr	6820	26656
x"00",	-- Hex Addr	6821	26657
x"00",	-- Hex Addr	6822	26658
x"00",	-- Hex Addr	6823	26659
x"00",	-- Hex Addr	6824	26660
x"00",	-- Hex Addr	6825	26661
x"00",	-- Hex Addr	6826	26662
x"00",	-- Hex Addr	6827	26663
x"00",	-- Hex Addr	6828	26664
x"00",	-- Hex Addr	6829	26665
x"00",	-- Hex Addr	682A	26666
x"00",	-- Hex Addr	682B	26667
x"00",	-- Hex Addr	682C	26668
x"00",	-- Hex Addr	682D	26669
x"00",	-- Hex Addr	682E	26670
x"00",	-- Hex Addr	682F	26671
x"00",	-- Hex Addr	6830	26672
x"00",	-- Hex Addr	6831	26673
x"00",	-- Hex Addr	6832	26674
x"00",	-- Hex Addr	6833	26675
x"00",	-- Hex Addr	6834	26676
x"00",	-- Hex Addr	6835	26677
x"00",	-- Hex Addr	6836	26678
x"00",	-- Hex Addr	6837	26679
x"00",	-- Hex Addr	6838	26680
x"00",	-- Hex Addr	6839	26681
x"00",	-- Hex Addr	683A	26682
x"00",	-- Hex Addr	683B	26683
x"00",	-- Hex Addr	683C	26684
x"00",	-- Hex Addr	683D	26685
x"00",	-- Hex Addr	683E	26686
x"00",	-- Hex Addr	683F	26687
x"00",	-- Hex Addr	6840	26688
x"00",	-- Hex Addr	6841	26689
x"00",	-- Hex Addr	6842	26690
x"00",	-- Hex Addr	6843	26691
x"00",	-- Hex Addr	6844	26692
x"00",	-- Hex Addr	6845	26693
x"00",	-- Hex Addr	6846	26694
x"00",	-- Hex Addr	6847	26695
x"00",	-- Hex Addr	6848	26696
x"00",	-- Hex Addr	6849	26697
x"00",	-- Hex Addr	684A	26698
x"00",	-- Hex Addr	684B	26699
x"00",	-- Hex Addr	684C	26700
x"00",	-- Hex Addr	684D	26701
x"00",	-- Hex Addr	684E	26702
x"00",	-- Hex Addr	684F	26703
x"00",	-- Hex Addr	6850	26704
x"00",	-- Hex Addr	6851	26705
x"00",	-- Hex Addr	6852	26706
x"00",	-- Hex Addr	6853	26707
x"00",	-- Hex Addr	6854	26708
x"00",	-- Hex Addr	6855	26709
x"00",	-- Hex Addr	6856	26710
x"00",	-- Hex Addr	6857	26711
x"00",	-- Hex Addr	6858	26712
x"00",	-- Hex Addr	6859	26713
x"00",	-- Hex Addr	685A	26714
x"00",	-- Hex Addr	685B	26715
x"00",	-- Hex Addr	685C	26716
x"00",	-- Hex Addr	685D	26717
x"00",	-- Hex Addr	685E	26718
x"00",	-- Hex Addr	685F	26719
x"00",	-- Hex Addr	6860	26720
x"00",	-- Hex Addr	6861	26721
x"00",	-- Hex Addr	6862	26722
x"00",	-- Hex Addr	6863	26723
x"00",	-- Hex Addr	6864	26724
x"00",	-- Hex Addr	6865	26725
x"00",	-- Hex Addr	6866	26726
x"00",	-- Hex Addr	6867	26727
x"00",	-- Hex Addr	6868	26728
x"00",	-- Hex Addr	6869	26729
x"00",	-- Hex Addr	686A	26730
x"00",	-- Hex Addr	686B	26731
x"00",	-- Hex Addr	686C	26732
x"00",	-- Hex Addr	686D	26733
x"00",	-- Hex Addr	686E	26734
x"00",	-- Hex Addr	686F	26735
x"00",	-- Hex Addr	6870	26736
x"00",	-- Hex Addr	6871	26737
x"00",	-- Hex Addr	6872	26738
x"00",	-- Hex Addr	6873	26739
x"00",	-- Hex Addr	6874	26740
x"00",	-- Hex Addr	6875	26741
x"00",	-- Hex Addr	6876	26742
x"00",	-- Hex Addr	6877	26743
x"00",	-- Hex Addr	6878	26744
x"00",	-- Hex Addr	6879	26745
x"00",	-- Hex Addr	687A	26746
x"00",	-- Hex Addr	687B	26747
x"00",	-- Hex Addr	687C	26748
x"00",	-- Hex Addr	687D	26749
x"00",	-- Hex Addr	687E	26750
x"00",	-- Hex Addr	687F	26751
x"00",	-- Hex Addr	6880	26752
x"00",	-- Hex Addr	6881	26753
x"00",	-- Hex Addr	6882	26754
x"00",	-- Hex Addr	6883	26755
x"00",	-- Hex Addr	6884	26756
x"00",	-- Hex Addr	6885	26757
x"00",	-- Hex Addr	6886	26758
x"00",	-- Hex Addr	6887	26759
x"00",	-- Hex Addr	6888	26760
x"00",	-- Hex Addr	6889	26761
x"00",	-- Hex Addr	688A	26762
x"00",	-- Hex Addr	688B	26763
x"00",	-- Hex Addr	688C	26764
x"00",	-- Hex Addr	688D	26765
x"00",	-- Hex Addr	688E	26766
x"00",	-- Hex Addr	688F	26767
x"00",	-- Hex Addr	6890	26768
x"00",	-- Hex Addr	6891	26769
x"00",	-- Hex Addr	6892	26770
x"00",	-- Hex Addr	6893	26771
x"00",	-- Hex Addr	6894	26772
x"00",	-- Hex Addr	6895	26773
x"00",	-- Hex Addr	6896	26774
x"00",	-- Hex Addr	6897	26775
x"00",	-- Hex Addr	6898	26776
x"00",	-- Hex Addr	6899	26777
x"00",	-- Hex Addr	689A	26778
x"00",	-- Hex Addr	689B	26779
x"00",	-- Hex Addr	689C	26780
x"00",	-- Hex Addr	689D	26781
x"00",	-- Hex Addr	689E	26782
x"00",	-- Hex Addr	689F	26783
x"00",	-- Hex Addr	68A0	26784
x"00",	-- Hex Addr	68A1	26785
x"00",	-- Hex Addr	68A2	26786
x"00",	-- Hex Addr	68A3	26787
x"00",	-- Hex Addr	68A4	26788
x"00",	-- Hex Addr	68A5	26789
x"00",	-- Hex Addr	68A6	26790
x"00",	-- Hex Addr	68A7	26791
x"00",	-- Hex Addr	68A8	26792
x"00",	-- Hex Addr	68A9	26793
x"00",	-- Hex Addr	68AA	26794
x"00",	-- Hex Addr	68AB	26795
x"00",	-- Hex Addr	68AC	26796
x"00",	-- Hex Addr	68AD	26797
x"00",	-- Hex Addr	68AE	26798
x"00",	-- Hex Addr	68AF	26799
x"00",	-- Hex Addr	68B0	26800
x"00",	-- Hex Addr	68B1	26801
x"00",	-- Hex Addr	68B2	26802
x"00",	-- Hex Addr	68B3	26803
x"00",	-- Hex Addr	68B4	26804
x"00",	-- Hex Addr	68B5	26805
x"00",	-- Hex Addr	68B6	26806
x"00",	-- Hex Addr	68B7	26807
x"00",	-- Hex Addr	68B8	26808
x"00",	-- Hex Addr	68B9	26809
x"00",	-- Hex Addr	68BA	26810
x"00",	-- Hex Addr	68BB	26811
x"00",	-- Hex Addr	68BC	26812
x"00",	-- Hex Addr	68BD	26813
x"00",	-- Hex Addr	68BE	26814
x"00",	-- Hex Addr	68BF	26815
x"00",	-- Hex Addr	68C0	26816
x"00",	-- Hex Addr	68C1	26817
x"00",	-- Hex Addr	68C2	26818
x"00",	-- Hex Addr	68C3	26819
x"00",	-- Hex Addr	68C4	26820
x"00",	-- Hex Addr	68C5	26821
x"00",	-- Hex Addr	68C6	26822
x"00",	-- Hex Addr	68C7	26823
x"00",	-- Hex Addr	68C8	26824
x"00",	-- Hex Addr	68C9	26825
x"00",	-- Hex Addr	68CA	26826
x"00",	-- Hex Addr	68CB	26827
x"00",	-- Hex Addr	68CC	26828
x"00",	-- Hex Addr	68CD	26829
x"00",	-- Hex Addr	68CE	26830
x"00",	-- Hex Addr	68CF	26831
x"00",	-- Hex Addr	68D0	26832
x"00",	-- Hex Addr	68D1	26833
x"00",	-- Hex Addr	68D2	26834
x"00",	-- Hex Addr	68D3	26835
x"00",	-- Hex Addr	68D4	26836
x"00",	-- Hex Addr	68D5	26837
x"00",	-- Hex Addr	68D6	26838
x"00",	-- Hex Addr	68D7	26839
x"00",	-- Hex Addr	68D8	26840
x"00",	-- Hex Addr	68D9	26841
x"00",	-- Hex Addr	68DA	26842
x"00",	-- Hex Addr	68DB	26843
x"00",	-- Hex Addr	68DC	26844
x"00",	-- Hex Addr	68DD	26845
x"00",	-- Hex Addr	68DE	26846
x"00",	-- Hex Addr	68DF	26847
x"00",	-- Hex Addr	68E0	26848
x"00",	-- Hex Addr	68E1	26849
x"00",	-- Hex Addr	68E2	26850
x"00",	-- Hex Addr	68E3	26851
x"00",	-- Hex Addr	68E4	26852
x"00",	-- Hex Addr	68E5	26853
x"00",	-- Hex Addr	68E6	26854
x"00",	-- Hex Addr	68E7	26855
x"00",	-- Hex Addr	68E8	26856
x"00",	-- Hex Addr	68E9	26857
x"00",	-- Hex Addr	68EA	26858
x"00",	-- Hex Addr	68EB	26859
x"00",	-- Hex Addr	68EC	26860
x"00",	-- Hex Addr	68ED	26861
x"00",	-- Hex Addr	68EE	26862
x"00",	-- Hex Addr	68EF	26863
x"00",	-- Hex Addr	68F0	26864
x"00",	-- Hex Addr	68F1	26865
x"00",	-- Hex Addr	68F2	26866
x"00",	-- Hex Addr	68F3	26867
x"00",	-- Hex Addr	68F4	26868
x"00",	-- Hex Addr	68F5	26869
x"00",	-- Hex Addr	68F6	26870
x"00",	-- Hex Addr	68F7	26871
x"00",	-- Hex Addr	68F8	26872
x"00",	-- Hex Addr	68F9	26873
x"00",	-- Hex Addr	68FA	26874
x"00",	-- Hex Addr	68FB	26875
x"00",	-- Hex Addr	68FC	26876
x"00",	-- Hex Addr	68FD	26877
x"00",	-- Hex Addr	68FE	26878
x"00",	-- Hex Addr	68FF	26879
x"00",	-- Hex Addr	6900	26880
x"00",	-- Hex Addr	6901	26881
x"00",	-- Hex Addr	6902	26882
x"00",	-- Hex Addr	6903	26883
x"00",	-- Hex Addr	6904	26884
x"00",	-- Hex Addr	6905	26885
x"00",	-- Hex Addr	6906	26886
x"00",	-- Hex Addr	6907	26887
x"00",	-- Hex Addr	6908	26888
x"00",	-- Hex Addr	6909	26889
x"00",	-- Hex Addr	690A	26890
x"00",	-- Hex Addr	690B	26891
x"00",	-- Hex Addr	690C	26892
x"00",	-- Hex Addr	690D	26893
x"00",	-- Hex Addr	690E	26894
x"00",	-- Hex Addr	690F	26895
x"00",	-- Hex Addr	6910	26896
x"00",	-- Hex Addr	6911	26897
x"00",	-- Hex Addr	6912	26898
x"00",	-- Hex Addr	6913	26899
x"00",	-- Hex Addr	6914	26900
x"00",	-- Hex Addr	6915	26901
x"00",	-- Hex Addr	6916	26902
x"00",	-- Hex Addr	6917	26903
x"00",	-- Hex Addr	6918	26904
x"00",	-- Hex Addr	6919	26905
x"00",	-- Hex Addr	691A	26906
x"00",	-- Hex Addr	691B	26907
x"00",	-- Hex Addr	691C	26908
x"00",	-- Hex Addr	691D	26909
x"00",	-- Hex Addr	691E	26910
x"00",	-- Hex Addr	691F	26911
x"00",	-- Hex Addr	6920	26912
x"00",	-- Hex Addr	6921	26913
x"00",	-- Hex Addr	6922	26914
x"00",	-- Hex Addr	6923	26915
x"00",	-- Hex Addr	6924	26916
x"00",	-- Hex Addr	6925	26917
x"00",	-- Hex Addr	6926	26918
x"00",	-- Hex Addr	6927	26919
x"00",	-- Hex Addr	6928	26920
x"00",	-- Hex Addr	6929	26921
x"00",	-- Hex Addr	692A	26922
x"00",	-- Hex Addr	692B	26923
x"00",	-- Hex Addr	692C	26924
x"00",	-- Hex Addr	692D	26925
x"00",	-- Hex Addr	692E	26926
x"00",	-- Hex Addr	692F	26927
x"00",	-- Hex Addr	6930	26928
x"00",	-- Hex Addr	6931	26929
x"00",	-- Hex Addr	6932	26930
x"00",	-- Hex Addr	6933	26931
x"00",	-- Hex Addr	6934	26932
x"00",	-- Hex Addr	6935	26933
x"00",	-- Hex Addr	6936	26934
x"00",	-- Hex Addr	6937	26935
x"00",	-- Hex Addr	6938	26936
x"00",	-- Hex Addr	6939	26937
x"00",	-- Hex Addr	693A	26938
x"00",	-- Hex Addr	693B	26939
x"00",	-- Hex Addr	693C	26940
x"00",	-- Hex Addr	693D	26941
x"00",	-- Hex Addr	693E	26942
x"00",	-- Hex Addr	693F	26943
x"00",	-- Hex Addr	6940	26944
x"00",	-- Hex Addr	6941	26945
x"00",	-- Hex Addr	6942	26946
x"00",	-- Hex Addr	6943	26947
x"00",	-- Hex Addr	6944	26948
x"00",	-- Hex Addr	6945	26949
x"00",	-- Hex Addr	6946	26950
x"00",	-- Hex Addr	6947	26951
x"00",	-- Hex Addr	6948	26952
x"00",	-- Hex Addr	6949	26953
x"00",	-- Hex Addr	694A	26954
x"00",	-- Hex Addr	694B	26955
x"00",	-- Hex Addr	694C	26956
x"00",	-- Hex Addr	694D	26957
x"00",	-- Hex Addr	694E	26958
x"00",	-- Hex Addr	694F	26959
x"00",	-- Hex Addr	6950	26960
x"00",	-- Hex Addr	6951	26961
x"00",	-- Hex Addr	6952	26962
x"00",	-- Hex Addr	6953	26963
x"00",	-- Hex Addr	6954	26964
x"00",	-- Hex Addr	6955	26965
x"00",	-- Hex Addr	6956	26966
x"00",	-- Hex Addr	6957	26967
x"00",	-- Hex Addr	6958	26968
x"00",	-- Hex Addr	6959	26969
x"00",	-- Hex Addr	695A	26970
x"00",	-- Hex Addr	695B	26971
x"00",	-- Hex Addr	695C	26972
x"00",	-- Hex Addr	695D	26973
x"00",	-- Hex Addr	695E	26974
x"00",	-- Hex Addr	695F	26975
x"00",	-- Hex Addr	6960	26976
x"00",	-- Hex Addr	6961	26977
x"00",	-- Hex Addr	6962	26978
x"00",	-- Hex Addr	6963	26979
x"00",	-- Hex Addr	6964	26980
x"00",	-- Hex Addr	6965	26981
x"00",	-- Hex Addr	6966	26982
x"00",	-- Hex Addr	6967	26983
x"00",	-- Hex Addr	6968	26984
x"00",	-- Hex Addr	6969	26985
x"00",	-- Hex Addr	696A	26986
x"00",	-- Hex Addr	696B	26987
x"00",	-- Hex Addr	696C	26988
x"00",	-- Hex Addr	696D	26989
x"00",	-- Hex Addr	696E	26990
x"00",	-- Hex Addr	696F	26991
x"00",	-- Hex Addr	6970	26992
x"00",	-- Hex Addr	6971	26993
x"00",	-- Hex Addr	6972	26994
x"00",	-- Hex Addr	6973	26995
x"00",	-- Hex Addr	6974	26996
x"00",	-- Hex Addr	6975	26997
x"00",	-- Hex Addr	6976	26998
x"00",	-- Hex Addr	6977	26999
x"00",	-- Hex Addr	6978	27000
x"00",	-- Hex Addr	6979	27001
x"00",	-- Hex Addr	697A	27002
x"00",	-- Hex Addr	697B	27003
x"00",	-- Hex Addr	697C	27004
x"00",	-- Hex Addr	697D	27005
x"00",	-- Hex Addr	697E	27006
x"00",	-- Hex Addr	697F	27007
x"00",	-- Hex Addr	6980	27008
x"00",	-- Hex Addr	6981	27009
x"00",	-- Hex Addr	6982	27010
x"00",	-- Hex Addr	6983	27011
x"00",	-- Hex Addr	6984	27012
x"00",	-- Hex Addr	6985	27013
x"00",	-- Hex Addr	6986	27014
x"00",	-- Hex Addr	6987	27015
x"00",	-- Hex Addr	6988	27016
x"00",	-- Hex Addr	6989	27017
x"00",	-- Hex Addr	698A	27018
x"00",	-- Hex Addr	698B	27019
x"00",	-- Hex Addr	698C	27020
x"00",	-- Hex Addr	698D	27021
x"00",	-- Hex Addr	698E	27022
x"00",	-- Hex Addr	698F	27023
x"00",	-- Hex Addr	6990	27024
x"00",	-- Hex Addr	6991	27025
x"00",	-- Hex Addr	6992	27026
x"00",	-- Hex Addr	6993	27027
x"00",	-- Hex Addr	6994	27028
x"00",	-- Hex Addr	6995	27029
x"00",	-- Hex Addr	6996	27030
x"00",	-- Hex Addr	6997	27031
x"00",	-- Hex Addr	6998	27032
x"00",	-- Hex Addr	6999	27033
x"00",	-- Hex Addr	699A	27034
x"00",	-- Hex Addr	699B	27035
x"00",	-- Hex Addr	699C	27036
x"00",	-- Hex Addr	699D	27037
x"00",	-- Hex Addr	699E	27038
x"00",	-- Hex Addr	699F	27039
x"00",	-- Hex Addr	69A0	27040
x"00",	-- Hex Addr	69A1	27041
x"00",	-- Hex Addr	69A2	27042
x"00",	-- Hex Addr	69A3	27043
x"00",	-- Hex Addr	69A4	27044
x"00",	-- Hex Addr	69A5	27045
x"00",	-- Hex Addr	69A6	27046
x"00",	-- Hex Addr	69A7	27047
x"00",	-- Hex Addr	69A8	27048
x"00",	-- Hex Addr	69A9	27049
x"00",	-- Hex Addr	69AA	27050
x"00",	-- Hex Addr	69AB	27051
x"00",	-- Hex Addr	69AC	27052
x"00",	-- Hex Addr	69AD	27053
x"00",	-- Hex Addr	69AE	27054
x"00",	-- Hex Addr	69AF	27055
x"00",	-- Hex Addr	69B0	27056
x"00",	-- Hex Addr	69B1	27057
x"00",	-- Hex Addr	69B2	27058
x"00",	-- Hex Addr	69B3	27059
x"00",	-- Hex Addr	69B4	27060
x"00",	-- Hex Addr	69B5	27061
x"00",	-- Hex Addr	69B6	27062
x"00",	-- Hex Addr	69B7	27063
x"00",	-- Hex Addr	69B8	27064
x"00",	-- Hex Addr	69B9	27065
x"00",	-- Hex Addr	69BA	27066
x"00",	-- Hex Addr	69BB	27067
x"00",	-- Hex Addr	69BC	27068
x"00",	-- Hex Addr	69BD	27069
x"00",	-- Hex Addr	69BE	27070
x"00",	-- Hex Addr	69BF	27071
x"00",	-- Hex Addr	69C0	27072
x"00",	-- Hex Addr	69C1	27073
x"00",	-- Hex Addr	69C2	27074
x"00",	-- Hex Addr	69C3	27075
x"00",	-- Hex Addr	69C4	27076
x"00",	-- Hex Addr	69C5	27077
x"00",	-- Hex Addr	69C6	27078
x"00",	-- Hex Addr	69C7	27079
x"00",	-- Hex Addr	69C8	27080
x"00",	-- Hex Addr	69C9	27081
x"00",	-- Hex Addr	69CA	27082
x"00",	-- Hex Addr	69CB	27083
x"00",	-- Hex Addr	69CC	27084
x"00",	-- Hex Addr	69CD	27085
x"00",	-- Hex Addr	69CE	27086
x"00",	-- Hex Addr	69CF	27087
x"00",	-- Hex Addr	69D0	27088
x"00",	-- Hex Addr	69D1	27089
x"00",	-- Hex Addr	69D2	27090
x"00",	-- Hex Addr	69D3	27091
x"00",	-- Hex Addr	69D4	27092
x"00",	-- Hex Addr	69D5	27093
x"00",	-- Hex Addr	69D6	27094
x"00",	-- Hex Addr	69D7	27095
x"00",	-- Hex Addr	69D8	27096
x"00",	-- Hex Addr	69D9	27097
x"00",	-- Hex Addr	69DA	27098
x"00",	-- Hex Addr	69DB	27099
x"00",	-- Hex Addr	69DC	27100
x"00",	-- Hex Addr	69DD	27101
x"00",	-- Hex Addr	69DE	27102
x"00",	-- Hex Addr	69DF	27103
x"00",	-- Hex Addr	69E0	27104
x"00",	-- Hex Addr	69E1	27105
x"00",	-- Hex Addr	69E2	27106
x"00",	-- Hex Addr	69E3	27107
x"00",	-- Hex Addr	69E4	27108
x"00",	-- Hex Addr	69E5	27109
x"00",	-- Hex Addr	69E6	27110
x"00",	-- Hex Addr	69E7	27111
x"00",	-- Hex Addr	69E8	27112
x"00",	-- Hex Addr	69E9	27113
x"00",	-- Hex Addr	69EA	27114
x"00",	-- Hex Addr	69EB	27115
x"00",	-- Hex Addr	69EC	27116
x"00",	-- Hex Addr	69ED	27117
x"00",	-- Hex Addr	69EE	27118
x"00",	-- Hex Addr	69EF	27119
x"00",	-- Hex Addr	69F0	27120
x"00",	-- Hex Addr	69F1	27121
x"00",	-- Hex Addr	69F2	27122
x"00",	-- Hex Addr	69F3	27123
x"00",	-- Hex Addr	69F4	27124
x"00",	-- Hex Addr	69F5	27125
x"00",	-- Hex Addr	69F6	27126
x"00",	-- Hex Addr	69F7	27127
x"00",	-- Hex Addr	69F8	27128
x"00",	-- Hex Addr	69F9	27129
x"00",	-- Hex Addr	69FA	27130
x"00",	-- Hex Addr	69FB	27131
x"00",	-- Hex Addr	69FC	27132
x"00",	-- Hex Addr	69FD	27133
x"00",	-- Hex Addr	69FE	27134
x"00",	-- Hex Addr	69FF	27135
x"00",	-- Hex Addr	6A00	27136
x"00",	-- Hex Addr	6A01	27137
x"00",	-- Hex Addr	6A02	27138
x"00",	-- Hex Addr	6A03	27139
x"00",	-- Hex Addr	6A04	27140
x"00",	-- Hex Addr	6A05	27141
x"00",	-- Hex Addr	6A06	27142
x"00",	-- Hex Addr	6A07	27143
x"00",	-- Hex Addr	6A08	27144
x"00",	-- Hex Addr	6A09	27145
x"00",	-- Hex Addr	6A0A	27146
x"00",	-- Hex Addr	6A0B	27147
x"00",	-- Hex Addr	6A0C	27148
x"00",	-- Hex Addr	6A0D	27149
x"00",	-- Hex Addr	6A0E	27150
x"00",	-- Hex Addr	6A0F	27151
x"00",	-- Hex Addr	6A10	27152
x"00",	-- Hex Addr	6A11	27153
x"00",	-- Hex Addr	6A12	27154
x"00",	-- Hex Addr	6A13	27155
x"00",	-- Hex Addr	6A14	27156
x"00",	-- Hex Addr	6A15	27157
x"00",	-- Hex Addr	6A16	27158
x"00",	-- Hex Addr	6A17	27159
x"00",	-- Hex Addr	6A18	27160
x"00",	-- Hex Addr	6A19	27161
x"00",	-- Hex Addr	6A1A	27162
x"00",	-- Hex Addr	6A1B	27163
x"00",	-- Hex Addr	6A1C	27164
x"00",	-- Hex Addr	6A1D	27165
x"00",	-- Hex Addr	6A1E	27166
x"00",	-- Hex Addr	6A1F	27167
x"00",	-- Hex Addr	6A20	27168
x"00",	-- Hex Addr	6A21	27169
x"00",	-- Hex Addr	6A22	27170
x"00",	-- Hex Addr	6A23	27171
x"00",	-- Hex Addr	6A24	27172
x"00",	-- Hex Addr	6A25	27173
x"00",	-- Hex Addr	6A26	27174
x"00",	-- Hex Addr	6A27	27175
x"00",	-- Hex Addr	6A28	27176
x"00",	-- Hex Addr	6A29	27177
x"00",	-- Hex Addr	6A2A	27178
x"00",	-- Hex Addr	6A2B	27179
x"00",	-- Hex Addr	6A2C	27180
x"00",	-- Hex Addr	6A2D	27181
x"00",	-- Hex Addr	6A2E	27182
x"00",	-- Hex Addr	6A2F	27183
x"00",	-- Hex Addr	6A30	27184
x"00",	-- Hex Addr	6A31	27185
x"00",	-- Hex Addr	6A32	27186
x"00",	-- Hex Addr	6A33	27187
x"00",	-- Hex Addr	6A34	27188
x"00",	-- Hex Addr	6A35	27189
x"00",	-- Hex Addr	6A36	27190
x"00",	-- Hex Addr	6A37	27191
x"00",	-- Hex Addr	6A38	27192
x"00",	-- Hex Addr	6A39	27193
x"00",	-- Hex Addr	6A3A	27194
x"00",	-- Hex Addr	6A3B	27195
x"00",	-- Hex Addr	6A3C	27196
x"00",	-- Hex Addr	6A3D	27197
x"00",	-- Hex Addr	6A3E	27198
x"00",	-- Hex Addr	6A3F	27199
x"00",	-- Hex Addr	6A40	27200
x"00",	-- Hex Addr	6A41	27201
x"00",	-- Hex Addr	6A42	27202
x"00",	-- Hex Addr	6A43	27203
x"00",	-- Hex Addr	6A44	27204
x"00",	-- Hex Addr	6A45	27205
x"00",	-- Hex Addr	6A46	27206
x"00",	-- Hex Addr	6A47	27207
x"00",	-- Hex Addr	6A48	27208
x"00",	-- Hex Addr	6A49	27209
x"00",	-- Hex Addr	6A4A	27210
x"00",	-- Hex Addr	6A4B	27211
x"00",	-- Hex Addr	6A4C	27212
x"00",	-- Hex Addr	6A4D	27213
x"00",	-- Hex Addr	6A4E	27214
x"00",	-- Hex Addr	6A4F	27215
x"00",	-- Hex Addr	6A50	27216
x"00",	-- Hex Addr	6A51	27217
x"00",	-- Hex Addr	6A52	27218
x"00",	-- Hex Addr	6A53	27219
x"00",	-- Hex Addr	6A54	27220
x"00",	-- Hex Addr	6A55	27221
x"00",	-- Hex Addr	6A56	27222
x"00",	-- Hex Addr	6A57	27223
x"00",	-- Hex Addr	6A58	27224
x"00",	-- Hex Addr	6A59	27225
x"00",	-- Hex Addr	6A5A	27226
x"00",	-- Hex Addr	6A5B	27227
x"00",	-- Hex Addr	6A5C	27228
x"00",	-- Hex Addr	6A5D	27229
x"00",	-- Hex Addr	6A5E	27230
x"00",	-- Hex Addr	6A5F	27231
x"00",	-- Hex Addr	6A60	27232
x"00",	-- Hex Addr	6A61	27233
x"00",	-- Hex Addr	6A62	27234
x"00",	-- Hex Addr	6A63	27235
x"00",	-- Hex Addr	6A64	27236
x"00",	-- Hex Addr	6A65	27237
x"00",	-- Hex Addr	6A66	27238
x"00",	-- Hex Addr	6A67	27239
x"00",	-- Hex Addr	6A68	27240
x"00",	-- Hex Addr	6A69	27241
x"00",	-- Hex Addr	6A6A	27242
x"00",	-- Hex Addr	6A6B	27243
x"00",	-- Hex Addr	6A6C	27244
x"00",	-- Hex Addr	6A6D	27245
x"00",	-- Hex Addr	6A6E	27246
x"00",	-- Hex Addr	6A6F	27247
x"00",	-- Hex Addr	6A70	27248
x"00",	-- Hex Addr	6A71	27249
x"00",	-- Hex Addr	6A72	27250
x"00",	-- Hex Addr	6A73	27251
x"00",	-- Hex Addr	6A74	27252
x"00",	-- Hex Addr	6A75	27253
x"00",	-- Hex Addr	6A76	27254
x"00",	-- Hex Addr	6A77	27255
x"00",	-- Hex Addr	6A78	27256
x"00",	-- Hex Addr	6A79	27257
x"00",	-- Hex Addr	6A7A	27258
x"00",	-- Hex Addr	6A7B	27259
x"00",	-- Hex Addr	6A7C	27260
x"00",	-- Hex Addr	6A7D	27261
x"00",	-- Hex Addr	6A7E	27262
x"00",	-- Hex Addr	6A7F	27263
x"00",	-- Hex Addr	6A80	27264
x"00",	-- Hex Addr	6A81	27265
x"00",	-- Hex Addr	6A82	27266
x"00",	-- Hex Addr	6A83	27267
x"00",	-- Hex Addr	6A84	27268
x"00",	-- Hex Addr	6A85	27269
x"00",	-- Hex Addr	6A86	27270
x"00",	-- Hex Addr	6A87	27271
x"00",	-- Hex Addr	6A88	27272
x"00",	-- Hex Addr	6A89	27273
x"00",	-- Hex Addr	6A8A	27274
x"00",	-- Hex Addr	6A8B	27275
x"00",	-- Hex Addr	6A8C	27276
x"00",	-- Hex Addr	6A8D	27277
x"00",	-- Hex Addr	6A8E	27278
x"00",	-- Hex Addr	6A8F	27279
x"00",	-- Hex Addr	6A90	27280
x"00",	-- Hex Addr	6A91	27281
x"00",	-- Hex Addr	6A92	27282
x"00",	-- Hex Addr	6A93	27283
x"00",	-- Hex Addr	6A94	27284
x"00",	-- Hex Addr	6A95	27285
x"00",	-- Hex Addr	6A96	27286
x"00",	-- Hex Addr	6A97	27287
x"00",	-- Hex Addr	6A98	27288
x"00",	-- Hex Addr	6A99	27289
x"00",	-- Hex Addr	6A9A	27290
x"00",	-- Hex Addr	6A9B	27291
x"00",	-- Hex Addr	6A9C	27292
x"00",	-- Hex Addr	6A9D	27293
x"00",	-- Hex Addr	6A9E	27294
x"00",	-- Hex Addr	6A9F	27295
x"00",	-- Hex Addr	6AA0	27296
x"00",	-- Hex Addr	6AA1	27297
x"00",	-- Hex Addr	6AA2	27298
x"00",	-- Hex Addr	6AA3	27299
x"00",	-- Hex Addr	6AA4	27300
x"00",	-- Hex Addr	6AA5	27301
x"00",	-- Hex Addr	6AA6	27302
x"00",	-- Hex Addr	6AA7	27303
x"00",	-- Hex Addr	6AA8	27304
x"00",	-- Hex Addr	6AA9	27305
x"00",	-- Hex Addr	6AAA	27306
x"00",	-- Hex Addr	6AAB	27307
x"00",	-- Hex Addr	6AAC	27308
x"00",	-- Hex Addr	6AAD	27309
x"00",	-- Hex Addr	6AAE	27310
x"00",	-- Hex Addr	6AAF	27311
x"00",	-- Hex Addr	6AB0	27312
x"00",	-- Hex Addr	6AB1	27313
x"00",	-- Hex Addr	6AB2	27314
x"00",	-- Hex Addr	6AB3	27315
x"00",	-- Hex Addr	6AB4	27316
x"00",	-- Hex Addr	6AB5	27317
x"00",	-- Hex Addr	6AB6	27318
x"00",	-- Hex Addr	6AB7	27319
x"00",	-- Hex Addr	6AB8	27320
x"00",	-- Hex Addr	6AB9	27321
x"00",	-- Hex Addr	6ABA	27322
x"00",	-- Hex Addr	6ABB	27323
x"00",	-- Hex Addr	6ABC	27324
x"00",	-- Hex Addr	6ABD	27325
x"00",	-- Hex Addr	6ABE	27326
x"00",	-- Hex Addr	6ABF	27327
x"00",	-- Hex Addr	6AC0	27328
x"00",	-- Hex Addr	6AC1	27329
x"00",	-- Hex Addr	6AC2	27330
x"00",	-- Hex Addr	6AC3	27331
x"00",	-- Hex Addr	6AC4	27332
x"00",	-- Hex Addr	6AC5	27333
x"00",	-- Hex Addr	6AC6	27334
x"00",	-- Hex Addr	6AC7	27335
x"00",	-- Hex Addr	6AC8	27336
x"00",	-- Hex Addr	6AC9	27337
x"00",	-- Hex Addr	6ACA	27338
x"00",	-- Hex Addr	6ACB	27339
x"00",	-- Hex Addr	6ACC	27340
x"00",	-- Hex Addr	6ACD	27341
x"00",	-- Hex Addr	6ACE	27342
x"00",	-- Hex Addr	6ACF	27343
x"00",	-- Hex Addr	6AD0	27344
x"00",	-- Hex Addr	6AD1	27345
x"00",	-- Hex Addr	6AD2	27346
x"00",	-- Hex Addr	6AD3	27347
x"00",	-- Hex Addr	6AD4	27348
x"00",	-- Hex Addr	6AD5	27349
x"00",	-- Hex Addr	6AD6	27350
x"00",	-- Hex Addr	6AD7	27351
x"00",	-- Hex Addr	6AD8	27352
x"00",	-- Hex Addr	6AD9	27353
x"00",	-- Hex Addr	6ADA	27354
x"00",	-- Hex Addr	6ADB	27355
x"00",	-- Hex Addr	6ADC	27356
x"00",	-- Hex Addr	6ADD	27357
x"00",	-- Hex Addr	6ADE	27358
x"00",	-- Hex Addr	6ADF	27359
x"00",	-- Hex Addr	6AE0	27360
x"00",	-- Hex Addr	6AE1	27361
x"00",	-- Hex Addr	6AE2	27362
x"00",	-- Hex Addr	6AE3	27363
x"00",	-- Hex Addr	6AE4	27364
x"00",	-- Hex Addr	6AE5	27365
x"00",	-- Hex Addr	6AE6	27366
x"00",	-- Hex Addr	6AE7	27367
x"00",	-- Hex Addr	6AE8	27368
x"00",	-- Hex Addr	6AE9	27369
x"00",	-- Hex Addr	6AEA	27370
x"00",	-- Hex Addr	6AEB	27371
x"00",	-- Hex Addr	6AEC	27372
x"00",	-- Hex Addr	6AED	27373
x"00",	-- Hex Addr	6AEE	27374
x"00",	-- Hex Addr	6AEF	27375
x"00",	-- Hex Addr	6AF0	27376
x"00",	-- Hex Addr	6AF1	27377
x"00",	-- Hex Addr	6AF2	27378
x"00",	-- Hex Addr	6AF3	27379
x"00",	-- Hex Addr	6AF4	27380
x"00",	-- Hex Addr	6AF5	27381
x"00",	-- Hex Addr	6AF6	27382
x"00",	-- Hex Addr	6AF7	27383
x"00",	-- Hex Addr	6AF8	27384
x"00",	-- Hex Addr	6AF9	27385
x"00",	-- Hex Addr	6AFA	27386
x"00",	-- Hex Addr	6AFB	27387
x"00",	-- Hex Addr	6AFC	27388
x"00",	-- Hex Addr	6AFD	27389
x"00",	-- Hex Addr	6AFE	27390
x"00",	-- Hex Addr	6AFF	27391
x"00",	-- Hex Addr	6B00	27392
x"00",	-- Hex Addr	6B01	27393
x"00",	-- Hex Addr	6B02	27394
x"00",	-- Hex Addr	6B03	27395
x"00",	-- Hex Addr	6B04	27396
x"00",	-- Hex Addr	6B05	27397
x"00",	-- Hex Addr	6B06	27398
x"00",	-- Hex Addr	6B07	27399
x"00",	-- Hex Addr	6B08	27400
x"00",	-- Hex Addr	6B09	27401
x"00",	-- Hex Addr	6B0A	27402
x"00",	-- Hex Addr	6B0B	27403
x"00",	-- Hex Addr	6B0C	27404
x"00",	-- Hex Addr	6B0D	27405
x"00",	-- Hex Addr	6B0E	27406
x"00",	-- Hex Addr	6B0F	27407
x"00",	-- Hex Addr	6B10	27408
x"00",	-- Hex Addr	6B11	27409
x"00",	-- Hex Addr	6B12	27410
x"00",	-- Hex Addr	6B13	27411
x"00",	-- Hex Addr	6B14	27412
x"00",	-- Hex Addr	6B15	27413
x"00",	-- Hex Addr	6B16	27414
x"00",	-- Hex Addr	6B17	27415
x"00",	-- Hex Addr	6B18	27416
x"00",	-- Hex Addr	6B19	27417
x"00",	-- Hex Addr	6B1A	27418
x"00",	-- Hex Addr	6B1B	27419
x"00",	-- Hex Addr	6B1C	27420
x"00",	-- Hex Addr	6B1D	27421
x"00",	-- Hex Addr	6B1E	27422
x"00",	-- Hex Addr	6B1F	27423
x"00",	-- Hex Addr	6B20	27424
x"00",	-- Hex Addr	6B21	27425
x"00",	-- Hex Addr	6B22	27426
x"00",	-- Hex Addr	6B23	27427
x"00",	-- Hex Addr	6B24	27428
x"00",	-- Hex Addr	6B25	27429
x"00",	-- Hex Addr	6B26	27430
x"00",	-- Hex Addr	6B27	27431
x"00",	-- Hex Addr	6B28	27432
x"00",	-- Hex Addr	6B29	27433
x"00",	-- Hex Addr	6B2A	27434
x"00",	-- Hex Addr	6B2B	27435
x"00",	-- Hex Addr	6B2C	27436
x"00",	-- Hex Addr	6B2D	27437
x"00",	-- Hex Addr	6B2E	27438
x"00",	-- Hex Addr	6B2F	27439
x"00",	-- Hex Addr	6B30	27440
x"00",	-- Hex Addr	6B31	27441
x"00",	-- Hex Addr	6B32	27442
x"00",	-- Hex Addr	6B33	27443
x"00",	-- Hex Addr	6B34	27444
x"00",	-- Hex Addr	6B35	27445
x"00",	-- Hex Addr	6B36	27446
x"00",	-- Hex Addr	6B37	27447
x"00",	-- Hex Addr	6B38	27448
x"00",	-- Hex Addr	6B39	27449
x"00",	-- Hex Addr	6B3A	27450
x"00",	-- Hex Addr	6B3B	27451
x"00",	-- Hex Addr	6B3C	27452
x"00",	-- Hex Addr	6B3D	27453
x"00",	-- Hex Addr	6B3E	27454
x"00",	-- Hex Addr	6B3F	27455
x"00",	-- Hex Addr	6B40	27456
x"00",	-- Hex Addr	6B41	27457
x"00",	-- Hex Addr	6B42	27458
x"00",	-- Hex Addr	6B43	27459
x"00",	-- Hex Addr	6B44	27460
x"00",	-- Hex Addr	6B45	27461
x"00",	-- Hex Addr	6B46	27462
x"00",	-- Hex Addr	6B47	27463
x"00",	-- Hex Addr	6B48	27464
x"00",	-- Hex Addr	6B49	27465
x"00",	-- Hex Addr	6B4A	27466
x"00",	-- Hex Addr	6B4B	27467
x"00",	-- Hex Addr	6B4C	27468
x"00",	-- Hex Addr	6B4D	27469
x"00",	-- Hex Addr	6B4E	27470
x"00",	-- Hex Addr	6B4F	27471
x"00",	-- Hex Addr	6B50	27472
x"00",	-- Hex Addr	6B51	27473
x"00",	-- Hex Addr	6B52	27474
x"00",	-- Hex Addr	6B53	27475
x"00",	-- Hex Addr	6B54	27476
x"00",	-- Hex Addr	6B55	27477
x"00",	-- Hex Addr	6B56	27478
x"00",	-- Hex Addr	6B57	27479
x"00",	-- Hex Addr	6B58	27480
x"00",	-- Hex Addr	6B59	27481
x"00",	-- Hex Addr	6B5A	27482
x"00",	-- Hex Addr	6B5B	27483
x"00",	-- Hex Addr	6B5C	27484
x"00",	-- Hex Addr	6B5D	27485
x"00",	-- Hex Addr	6B5E	27486
x"00",	-- Hex Addr	6B5F	27487
x"00",	-- Hex Addr	6B60	27488
x"00",	-- Hex Addr	6B61	27489
x"00",	-- Hex Addr	6B62	27490
x"00",	-- Hex Addr	6B63	27491
x"00",	-- Hex Addr	6B64	27492
x"00",	-- Hex Addr	6B65	27493
x"00",	-- Hex Addr	6B66	27494
x"00",	-- Hex Addr	6B67	27495
x"00",	-- Hex Addr	6B68	27496
x"00",	-- Hex Addr	6B69	27497
x"00",	-- Hex Addr	6B6A	27498
x"00",	-- Hex Addr	6B6B	27499
x"00",	-- Hex Addr	6B6C	27500
x"00",	-- Hex Addr	6B6D	27501
x"00",	-- Hex Addr	6B6E	27502
x"00",	-- Hex Addr	6B6F	27503
x"00",	-- Hex Addr	6B70	27504
x"00",	-- Hex Addr	6B71	27505
x"00",	-- Hex Addr	6B72	27506
x"00",	-- Hex Addr	6B73	27507
x"00",	-- Hex Addr	6B74	27508
x"00",	-- Hex Addr	6B75	27509
x"00",	-- Hex Addr	6B76	27510
x"00",	-- Hex Addr	6B77	27511
x"00",	-- Hex Addr	6B78	27512
x"00",	-- Hex Addr	6B79	27513
x"00",	-- Hex Addr	6B7A	27514
x"00",	-- Hex Addr	6B7B	27515
x"00",	-- Hex Addr	6B7C	27516
x"00",	-- Hex Addr	6B7D	27517
x"00",	-- Hex Addr	6B7E	27518
x"00",	-- Hex Addr	6B7F	27519
x"00",	-- Hex Addr	6B80	27520
x"00",	-- Hex Addr	6B81	27521
x"00",	-- Hex Addr	6B82	27522
x"00",	-- Hex Addr	6B83	27523
x"00",	-- Hex Addr	6B84	27524
x"00",	-- Hex Addr	6B85	27525
x"00",	-- Hex Addr	6B86	27526
x"00",	-- Hex Addr	6B87	27527
x"00",	-- Hex Addr	6B88	27528
x"00",	-- Hex Addr	6B89	27529
x"00",	-- Hex Addr	6B8A	27530
x"00",	-- Hex Addr	6B8B	27531
x"00",	-- Hex Addr	6B8C	27532
x"00",	-- Hex Addr	6B8D	27533
x"00",	-- Hex Addr	6B8E	27534
x"00",	-- Hex Addr	6B8F	27535
x"00",	-- Hex Addr	6B90	27536
x"00",	-- Hex Addr	6B91	27537
x"00",	-- Hex Addr	6B92	27538
x"00",	-- Hex Addr	6B93	27539
x"00",	-- Hex Addr	6B94	27540
x"00",	-- Hex Addr	6B95	27541
x"00",	-- Hex Addr	6B96	27542
x"00",	-- Hex Addr	6B97	27543
x"00",	-- Hex Addr	6B98	27544
x"00",	-- Hex Addr	6B99	27545
x"00",	-- Hex Addr	6B9A	27546
x"00",	-- Hex Addr	6B9B	27547
x"00",	-- Hex Addr	6B9C	27548
x"00",	-- Hex Addr	6B9D	27549
x"00",	-- Hex Addr	6B9E	27550
x"00",	-- Hex Addr	6B9F	27551
x"00",	-- Hex Addr	6BA0	27552
x"00",	-- Hex Addr	6BA1	27553
x"00",	-- Hex Addr	6BA2	27554
x"00",	-- Hex Addr	6BA3	27555
x"00",	-- Hex Addr	6BA4	27556
x"00",	-- Hex Addr	6BA5	27557
x"00",	-- Hex Addr	6BA6	27558
x"00",	-- Hex Addr	6BA7	27559
x"00",	-- Hex Addr	6BA8	27560
x"00",	-- Hex Addr	6BA9	27561
x"00",	-- Hex Addr	6BAA	27562
x"00",	-- Hex Addr	6BAB	27563
x"00",	-- Hex Addr	6BAC	27564
x"00",	-- Hex Addr	6BAD	27565
x"00",	-- Hex Addr	6BAE	27566
x"00",	-- Hex Addr	6BAF	27567
x"00",	-- Hex Addr	6BB0	27568
x"00",	-- Hex Addr	6BB1	27569
x"00",	-- Hex Addr	6BB2	27570
x"00",	-- Hex Addr	6BB3	27571
x"00",	-- Hex Addr	6BB4	27572
x"00",	-- Hex Addr	6BB5	27573
x"00",	-- Hex Addr	6BB6	27574
x"00",	-- Hex Addr	6BB7	27575
x"00",	-- Hex Addr	6BB8	27576
x"00",	-- Hex Addr	6BB9	27577
x"00",	-- Hex Addr	6BBA	27578
x"00",	-- Hex Addr	6BBB	27579
x"00",	-- Hex Addr	6BBC	27580
x"00",	-- Hex Addr	6BBD	27581
x"00",	-- Hex Addr	6BBE	27582
x"00",	-- Hex Addr	6BBF	27583
x"00",	-- Hex Addr	6BC0	27584
x"00",	-- Hex Addr	6BC1	27585
x"00",	-- Hex Addr	6BC2	27586
x"00",	-- Hex Addr	6BC3	27587
x"00",	-- Hex Addr	6BC4	27588
x"00",	-- Hex Addr	6BC5	27589
x"00",	-- Hex Addr	6BC6	27590
x"00",	-- Hex Addr	6BC7	27591
x"00",	-- Hex Addr	6BC8	27592
x"00",	-- Hex Addr	6BC9	27593
x"00",	-- Hex Addr	6BCA	27594
x"00",	-- Hex Addr	6BCB	27595
x"00",	-- Hex Addr	6BCC	27596
x"00",	-- Hex Addr	6BCD	27597
x"00",	-- Hex Addr	6BCE	27598
x"00",	-- Hex Addr	6BCF	27599
x"00",	-- Hex Addr	6BD0	27600
x"00",	-- Hex Addr	6BD1	27601
x"00",	-- Hex Addr	6BD2	27602
x"00",	-- Hex Addr	6BD3	27603
x"00",	-- Hex Addr	6BD4	27604
x"00",	-- Hex Addr	6BD5	27605
x"00",	-- Hex Addr	6BD6	27606
x"00",	-- Hex Addr	6BD7	27607
x"00",	-- Hex Addr	6BD8	27608
x"00",	-- Hex Addr	6BD9	27609
x"00",	-- Hex Addr	6BDA	27610
x"00",	-- Hex Addr	6BDB	27611
x"00",	-- Hex Addr	6BDC	27612
x"00",	-- Hex Addr	6BDD	27613
x"00",	-- Hex Addr	6BDE	27614
x"00",	-- Hex Addr	6BDF	27615
x"00",	-- Hex Addr	6BE0	27616
x"00",	-- Hex Addr	6BE1	27617
x"00",	-- Hex Addr	6BE2	27618
x"00",	-- Hex Addr	6BE3	27619
x"00",	-- Hex Addr	6BE4	27620
x"00",	-- Hex Addr	6BE5	27621
x"00",	-- Hex Addr	6BE6	27622
x"00",	-- Hex Addr	6BE7	27623
x"00",	-- Hex Addr	6BE8	27624
x"00",	-- Hex Addr	6BE9	27625
x"00",	-- Hex Addr	6BEA	27626
x"00",	-- Hex Addr	6BEB	27627
x"00",	-- Hex Addr	6BEC	27628
x"00",	-- Hex Addr	6BED	27629
x"00",	-- Hex Addr	6BEE	27630
x"00",	-- Hex Addr	6BEF	27631
x"00",	-- Hex Addr	6BF0	27632
x"00",	-- Hex Addr	6BF1	27633
x"00",	-- Hex Addr	6BF2	27634
x"00",	-- Hex Addr	6BF3	27635
x"00",	-- Hex Addr	6BF4	27636
x"00",	-- Hex Addr	6BF5	27637
x"00",	-- Hex Addr	6BF6	27638
x"00",	-- Hex Addr	6BF7	27639
x"00",	-- Hex Addr	6BF8	27640
x"00",	-- Hex Addr	6BF9	27641
x"00",	-- Hex Addr	6BFA	27642
x"00",	-- Hex Addr	6BFB	27643
x"00",	-- Hex Addr	6BFC	27644
x"00",	-- Hex Addr	6BFD	27645
x"00",	-- Hex Addr	6BFE	27646
x"00",	-- Hex Addr	6BFF	27647
x"00",	-- Hex Addr	6C00	27648
x"00",	-- Hex Addr	6C01	27649
x"00",	-- Hex Addr	6C02	27650
x"00",	-- Hex Addr	6C03	27651
x"00",	-- Hex Addr	6C04	27652
x"00",	-- Hex Addr	6C05	27653
x"00",	-- Hex Addr	6C06	27654
x"00",	-- Hex Addr	6C07	27655
x"00",	-- Hex Addr	6C08	27656
x"00",	-- Hex Addr	6C09	27657
x"00",	-- Hex Addr	6C0A	27658
x"00",	-- Hex Addr	6C0B	27659
x"00",	-- Hex Addr	6C0C	27660
x"00",	-- Hex Addr	6C0D	27661
x"00",	-- Hex Addr	6C0E	27662
x"00",	-- Hex Addr	6C0F	27663
x"00",	-- Hex Addr	6C10	27664
x"00",	-- Hex Addr	6C11	27665
x"00",	-- Hex Addr	6C12	27666
x"00",	-- Hex Addr	6C13	27667
x"00",	-- Hex Addr	6C14	27668
x"00",	-- Hex Addr	6C15	27669
x"00",	-- Hex Addr	6C16	27670
x"00",	-- Hex Addr	6C17	27671
x"00",	-- Hex Addr	6C18	27672
x"00",	-- Hex Addr	6C19	27673
x"00",	-- Hex Addr	6C1A	27674
x"00",	-- Hex Addr	6C1B	27675
x"00",	-- Hex Addr	6C1C	27676
x"00",	-- Hex Addr	6C1D	27677
x"00",	-- Hex Addr	6C1E	27678
x"00",	-- Hex Addr	6C1F	27679
x"00",	-- Hex Addr	6C20	27680
x"00",	-- Hex Addr	6C21	27681
x"00",	-- Hex Addr	6C22	27682
x"00",	-- Hex Addr	6C23	27683
x"00",	-- Hex Addr	6C24	27684
x"00",	-- Hex Addr	6C25	27685
x"00",	-- Hex Addr	6C26	27686
x"00",	-- Hex Addr	6C27	27687
x"00",	-- Hex Addr	6C28	27688
x"00",	-- Hex Addr	6C29	27689
x"00",	-- Hex Addr	6C2A	27690
x"00",	-- Hex Addr	6C2B	27691
x"00",	-- Hex Addr	6C2C	27692
x"00",	-- Hex Addr	6C2D	27693
x"00",	-- Hex Addr	6C2E	27694
x"00",	-- Hex Addr	6C2F	27695
x"00",	-- Hex Addr	6C30	27696
x"00",	-- Hex Addr	6C31	27697
x"00",	-- Hex Addr	6C32	27698
x"00",	-- Hex Addr	6C33	27699
x"00",	-- Hex Addr	6C34	27700
x"00",	-- Hex Addr	6C35	27701
x"00",	-- Hex Addr	6C36	27702
x"00",	-- Hex Addr	6C37	27703
x"00",	-- Hex Addr	6C38	27704
x"00",	-- Hex Addr	6C39	27705
x"00",	-- Hex Addr	6C3A	27706
x"00",	-- Hex Addr	6C3B	27707
x"00",	-- Hex Addr	6C3C	27708
x"00",	-- Hex Addr	6C3D	27709
x"00",	-- Hex Addr	6C3E	27710
x"00",	-- Hex Addr	6C3F	27711
x"00",	-- Hex Addr	6C40	27712
x"00",	-- Hex Addr	6C41	27713
x"00",	-- Hex Addr	6C42	27714
x"00",	-- Hex Addr	6C43	27715
x"00",	-- Hex Addr	6C44	27716
x"00",	-- Hex Addr	6C45	27717
x"00",	-- Hex Addr	6C46	27718
x"00",	-- Hex Addr	6C47	27719
x"00",	-- Hex Addr	6C48	27720
x"00",	-- Hex Addr	6C49	27721
x"00",	-- Hex Addr	6C4A	27722
x"00",	-- Hex Addr	6C4B	27723
x"00",	-- Hex Addr	6C4C	27724
x"00",	-- Hex Addr	6C4D	27725
x"00",	-- Hex Addr	6C4E	27726
x"00",	-- Hex Addr	6C4F	27727
x"00",	-- Hex Addr	6C50	27728
x"00",	-- Hex Addr	6C51	27729
x"00",	-- Hex Addr	6C52	27730
x"00",	-- Hex Addr	6C53	27731
x"00",	-- Hex Addr	6C54	27732
x"00",	-- Hex Addr	6C55	27733
x"00",	-- Hex Addr	6C56	27734
x"00",	-- Hex Addr	6C57	27735
x"00",	-- Hex Addr	6C58	27736
x"00",	-- Hex Addr	6C59	27737
x"00",	-- Hex Addr	6C5A	27738
x"00",	-- Hex Addr	6C5B	27739
x"00",	-- Hex Addr	6C5C	27740
x"00",	-- Hex Addr	6C5D	27741
x"00",	-- Hex Addr	6C5E	27742
x"00",	-- Hex Addr	6C5F	27743
x"00",	-- Hex Addr	6C60	27744
x"00",	-- Hex Addr	6C61	27745
x"00",	-- Hex Addr	6C62	27746
x"00",	-- Hex Addr	6C63	27747
x"00",	-- Hex Addr	6C64	27748
x"00",	-- Hex Addr	6C65	27749
x"00",	-- Hex Addr	6C66	27750
x"00",	-- Hex Addr	6C67	27751
x"00",	-- Hex Addr	6C68	27752
x"00",	-- Hex Addr	6C69	27753
x"00",	-- Hex Addr	6C6A	27754
x"00",	-- Hex Addr	6C6B	27755
x"00",	-- Hex Addr	6C6C	27756
x"00",	-- Hex Addr	6C6D	27757
x"00",	-- Hex Addr	6C6E	27758
x"00",	-- Hex Addr	6C6F	27759
x"00",	-- Hex Addr	6C70	27760
x"00",	-- Hex Addr	6C71	27761
x"00",	-- Hex Addr	6C72	27762
x"00",	-- Hex Addr	6C73	27763
x"00",	-- Hex Addr	6C74	27764
x"00",	-- Hex Addr	6C75	27765
x"00",	-- Hex Addr	6C76	27766
x"00",	-- Hex Addr	6C77	27767
x"00",	-- Hex Addr	6C78	27768
x"00",	-- Hex Addr	6C79	27769
x"00",	-- Hex Addr	6C7A	27770
x"00",	-- Hex Addr	6C7B	27771
x"00",	-- Hex Addr	6C7C	27772
x"00",	-- Hex Addr	6C7D	27773
x"00",	-- Hex Addr	6C7E	27774
x"00",	-- Hex Addr	6C7F	27775
x"00",	-- Hex Addr	6C80	27776
x"00",	-- Hex Addr	6C81	27777
x"00",	-- Hex Addr	6C82	27778
x"00",	-- Hex Addr	6C83	27779
x"00",	-- Hex Addr	6C84	27780
x"00",	-- Hex Addr	6C85	27781
x"00",	-- Hex Addr	6C86	27782
x"00",	-- Hex Addr	6C87	27783
x"00",	-- Hex Addr	6C88	27784
x"00",	-- Hex Addr	6C89	27785
x"00",	-- Hex Addr	6C8A	27786
x"00",	-- Hex Addr	6C8B	27787
x"00",	-- Hex Addr	6C8C	27788
x"00",	-- Hex Addr	6C8D	27789
x"00",	-- Hex Addr	6C8E	27790
x"00",	-- Hex Addr	6C8F	27791
x"00",	-- Hex Addr	6C90	27792
x"00",	-- Hex Addr	6C91	27793
x"00",	-- Hex Addr	6C92	27794
x"00",	-- Hex Addr	6C93	27795
x"00",	-- Hex Addr	6C94	27796
x"00",	-- Hex Addr	6C95	27797
x"00",	-- Hex Addr	6C96	27798
x"00",	-- Hex Addr	6C97	27799
x"00",	-- Hex Addr	6C98	27800
x"00",	-- Hex Addr	6C99	27801
x"00",	-- Hex Addr	6C9A	27802
x"00",	-- Hex Addr	6C9B	27803
x"00",	-- Hex Addr	6C9C	27804
x"00",	-- Hex Addr	6C9D	27805
x"00",	-- Hex Addr	6C9E	27806
x"00",	-- Hex Addr	6C9F	27807
x"00",	-- Hex Addr	6CA0	27808
x"00",	-- Hex Addr	6CA1	27809
x"00",	-- Hex Addr	6CA2	27810
x"00",	-- Hex Addr	6CA3	27811
x"00",	-- Hex Addr	6CA4	27812
x"00",	-- Hex Addr	6CA5	27813
x"00",	-- Hex Addr	6CA6	27814
x"00",	-- Hex Addr	6CA7	27815
x"00",	-- Hex Addr	6CA8	27816
x"00",	-- Hex Addr	6CA9	27817
x"00",	-- Hex Addr	6CAA	27818
x"00",	-- Hex Addr	6CAB	27819
x"00",	-- Hex Addr	6CAC	27820
x"00",	-- Hex Addr	6CAD	27821
x"00",	-- Hex Addr	6CAE	27822
x"00",	-- Hex Addr	6CAF	27823
x"00",	-- Hex Addr	6CB0	27824
x"00",	-- Hex Addr	6CB1	27825
x"00",	-- Hex Addr	6CB2	27826
x"00",	-- Hex Addr	6CB3	27827
x"00",	-- Hex Addr	6CB4	27828
x"00",	-- Hex Addr	6CB5	27829
x"00",	-- Hex Addr	6CB6	27830
x"00",	-- Hex Addr	6CB7	27831
x"00",	-- Hex Addr	6CB8	27832
x"00",	-- Hex Addr	6CB9	27833
x"00",	-- Hex Addr	6CBA	27834
x"00",	-- Hex Addr	6CBB	27835
x"00",	-- Hex Addr	6CBC	27836
x"00",	-- Hex Addr	6CBD	27837
x"00",	-- Hex Addr	6CBE	27838
x"00",	-- Hex Addr	6CBF	27839
x"00",	-- Hex Addr	6CC0	27840
x"00",	-- Hex Addr	6CC1	27841
x"00",	-- Hex Addr	6CC2	27842
x"00",	-- Hex Addr	6CC3	27843
x"00",	-- Hex Addr	6CC4	27844
x"00",	-- Hex Addr	6CC5	27845
x"00",	-- Hex Addr	6CC6	27846
x"00",	-- Hex Addr	6CC7	27847
x"00",	-- Hex Addr	6CC8	27848
x"00",	-- Hex Addr	6CC9	27849
x"00",	-- Hex Addr	6CCA	27850
x"00",	-- Hex Addr	6CCB	27851
x"00",	-- Hex Addr	6CCC	27852
x"00",	-- Hex Addr	6CCD	27853
x"00",	-- Hex Addr	6CCE	27854
x"00",	-- Hex Addr	6CCF	27855
x"00",	-- Hex Addr	6CD0	27856
x"00",	-- Hex Addr	6CD1	27857
x"00",	-- Hex Addr	6CD2	27858
x"00",	-- Hex Addr	6CD3	27859
x"00",	-- Hex Addr	6CD4	27860
x"00",	-- Hex Addr	6CD5	27861
x"00",	-- Hex Addr	6CD6	27862
x"00",	-- Hex Addr	6CD7	27863
x"00",	-- Hex Addr	6CD8	27864
x"00",	-- Hex Addr	6CD9	27865
x"00",	-- Hex Addr	6CDA	27866
x"00",	-- Hex Addr	6CDB	27867
x"00",	-- Hex Addr	6CDC	27868
x"00",	-- Hex Addr	6CDD	27869
x"00",	-- Hex Addr	6CDE	27870
x"00",	-- Hex Addr	6CDF	27871
x"00",	-- Hex Addr	6CE0	27872
x"00",	-- Hex Addr	6CE1	27873
x"00",	-- Hex Addr	6CE2	27874
x"00",	-- Hex Addr	6CE3	27875
x"00",	-- Hex Addr	6CE4	27876
x"00",	-- Hex Addr	6CE5	27877
x"00",	-- Hex Addr	6CE6	27878
x"00",	-- Hex Addr	6CE7	27879
x"00",	-- Hex Addr	6CE8	27880
x"00",	-- Hex Addr	6CE9	27881
x"00",	-- Hex Addr	6CEA	27882
x"00",	-- Hex Addr	6CEB	27883
x"00",	-- Hex Addr	6CEC	27884
x"00",	-- Hex Addr	6CED	27885
x"00",	-- Hex Addr	6CEE	27886
x"00",	-- Hex Addr	6CEF	27887
x"00",	-- Hex Addr	6CF0	27888
x"00",	-- Hex Addr	6CF1	27889
x"00",	-- Hex Addr	6CF2	27890
x"00",	-- Hex Addr	6CF3	27891
x"00",	-- Hex Addr	6CF4	27892
x"00",	-- Hex Addr	6CF5	27893
x"00",	-- Hex Addr	6CF6	27894
x"00",	-- Hex Addr	6CF7	27895
x"00",	-- Hex Addr	6CF8	27896
x"00",	-- Hex Addr	6CF9	27897
x"00",	-- Hex Addr	6CFA	27898
x"00",	-- Hex Addr	6CFB	27899
x"00",	-- Hex Addr	6CFC	27900
x"00",	-- Hex Addr	6CFD	27901
x"00",	-- Hex Addr	6CFE	27902
x"00",	-- Hex Addr	6CFF	27903
x"00",	-- Hex Addr	6D00	27904
x"00",	-- Hex Addr	6D01	27905
x"00",	-- Hex Addr	6D02	27906
x"00",	-- Hex Addr	6D03	27907
x"00",	-- Hex Addr	6D04	27908
x"00",	-- Hex Addr	6D05	27909
x"00",	-- Hex Addr	6D06	27910
x"00",	-- Hex Addr	6D07	27911
x"00",	-- Hex Addr	6D08	27912
x"00",	-- Hex Addr	6D09	27913
x"00",	-- Hex Addr	6D0A	27914
x"00",	-- Hex Addr	6D0B	27915
x"00",	-- Hex Addr	6D0C	27916
x"00",	-- Hex Addr	6D0D	27917
x"00",	-- Hex Addr	6D0E	27918
x"00",	-- Hex Addr	6D0F	27919
x"00",	-- Hex Addr	6D10	27920
x"00",	-- Hex Addr	6D11	27921
x"00",	-- Hex Addr	6D12	27922
x"00",	-- Hex Addr	6D13	27923
x"00",	-- Hex Addr	6D14	27924
x"00",	-- Hex Addr	6D15	27925
x"00",	-- Hex Addr	6D16	27926
x"00",	-- Hex Addr	6D17	27927
x"00",	-- Hex Addr	6D18	27928
x"00",	-- Hex Addr	6D19	27929
x"00",	-- Hex Addr	6D1A	27930
x"00",	-- Hex Addr	6D1B	27931
x"00",	-- Hex Addr	6D1C	27932
x"00",	-- Hex Addr	6D1D	27933
x"00",	-- Hex Addr	6D1E	27934
x"00",	-- Hex Addr	6D1F	27935
x"00",	-- Hex Addr	6D20	27936
x"00",	-- Hex Addr	6D21	27937
x"00",	-- Hex Addr	6D22	27938
x"00",	-- Hex Addr	6D23	27939
x"00",	-- Hex Addr	6D24	27940
x"00",	-- Hex Addr	6D25	27941
x"00",	-- Hex Addr	6D26	27942
x"00",	-- Hex Addr	6D27	27943
x"00",	-- Hex Addr	6D28	27944
x"00",	-- Hex Addr	6D29	27945
x"00",	-- Hex Addr	6D2A	27946
x"00",	-- Hex Addr	6D2B	27947
x"00",	-- Hex Addr	6D2C	27948
x"00",	-- Hex Addr	6D2D	27949
x"00",	-- Hex Addr	6D2E	27950
x"00",	-- Hex Addr	6D2F	27951
x"00",	-- Hex Addr	6D30	27952
x"00",	-- Hex Addr	6D31	27953
x"00",	-- Hex Addr	6D32	27954
x"00",	-- Hex Addr	6D33	27955
x"00",	-- Hex Addr	6D34	27956
x"00",	-- Hex Addr	6D35	27957
x"00",	-- Hex Addr	6D36	27958
x"00",	-- Hex Addr	6D37	27959
x"00",	-- Hex Addr	6D38	27960
x"00",	-- Hex Addr	6D39	27961
x"00",	-- Hex Addr	6D3A	27962
x"00",	-- Hex Addr	6D3B	27963
x"00",	-- Hex Addr	6D3C	27964
x"00",	-- Hex Addr	6D3D	27965
x"00",	-- Hex Addr	6D3E	27966
x"00",	-- Hex Addr	6D3F	27967
x"00",	-- Hex Addr	6D40	27968
x"00",	-- Hex Addr	6D41	27969
x"00",	-- Hex Addr	6D42	27970
x"00",	-- Hex Addr	6D43	27971
x"00",	-- Hex Addr	6D44	27972
x"00",	-- Hex Addr	6D45	27973
x"00",	-- Hex Addr	6D46	27974
x"00",	-- Hex Addr	6D47	27975
x"00",	-- Hex Addr	6D48	27976
x"00",	-- Hex Addr	6D49	27977
x"00",	-- Hex Addr	6D4A	27978
x"00",	-- Hex Addr	6D4B	27979
x"00",	-- Hex Addr	6D4C	27980
x"00",	-- Hex Addr	6D4D	27981
x"00",	-- Hex Addr	6D4E	27982
x"00",	-- Hex Addr	6D4F	27983
x"00",	-- Hex Addr	6D50	27984
x"00",	-- Hex Addr	6D51	27985
x"00",	-- Hex Addr	6D52	27986
x"00",	-- Hex Addr	6D53	27987
x"00",	-- Hex Addr	6D54	27988
x"00",	-- Hex Addr	6D55	27989
x"00",	-- Hex Addr	6D56	27990
x"00",	-- Hex Addr	6D57	27991
x"00",	-- Hex Addr	6D58	27992
x"00",	-- Hex Addr	6D59	27993
x"00",	-- Hex Addr	6D5A	27994
x"00",	-- Hex Addr	6D5B	27995
x"00",	-- Hex Addr	6D5C	27996
x"00",	-- Hex Addr	6D5D	27997
x"00",	-- Hex Addr	6D5E	27998
x"00",	-- Hex Addr	6D5F	27999
x"00",	-- Hex Addr	6D60	28000
x"00",	-- Hex Addr	6D61	28001
x"00",	-- Hex Addr	6D62	28002
x"00",	-- Hex Addr	6D63	28003
x"00",	-- Hex Addr	6D64	28004
x"00",	-- Hex Addr	6D65	28005
x"00",	-- Hex Addr	6D66	28006
x"00",	-- Hex Addr	6D67	28007
x"00",	-- Hex Addr	6D68	28008
x"00",	-- Hex Addr	6D69	28009
x"00",	-- Hex Addr	6D6A	28010
x"00",	-- Hex Addr	6D6B	28011
x"00",	-- Hex Addr	6D6C	28012
x"00",	-- Hex Addr	6D6D	28013
x"00",	-- Hex Addr	6D6E	28014
x"00",	-- Hex Addr	6D6F	28015
x"00",	-- Hex Addr	6D70	28016
x"00",	-- Hex Addr	6D71	28017
x"00",	-- Hex Addr	6D72	28018
x"00",	-- Hex Addr	6D73	28019
x"00",	-- Hex Addr	6D74	28020
x"00",	-- Hex Addr	6D75	28021
x"00",	-- Hex Addr	6D76	28022
x"00",	-- Hex Addr	6D77	28023
x"00",	-- Hex Addr	6D78	28024
x"00",	-- Hex Addr	6D79	28025
x"00",	-- Hex Addr	6D7A	28026
x"00",	-- Hex Addr	6D7B	28027
x"00",	-- Hex Addr	6D7C	28028
x"00",	-- Hex Addr	6D7D	28029
x"00",	-- Hex Addr	6D7E	28030
x"00",	-- Hex Addr	6D7F	28031
x"00",	-- Hex Addr	6D80	28032
x"00",	-- Hex Addr	6D81	28033
x"00",	-- Hex Addr	6D82	28034
x"00",	-- Hex Addr	6D83	28035
x"00",	-- Hex Addr	6D84	28036
x"00",	-- Hex Addr	6D85	28037
x"00",	-- Hex Addr	6D86	28038
x"00",	-- Hex Addr	6D87	28039
x"00",	-- Hex Addr	6D88	28040
x"00",	-- Hex Addr	6D89	28041
x"00",	-- Hex Addr	6D8A	28042
x"00",	-- Hex Addr	6D8B	28043
x"00",	-- Hex Addr	6D8C	28044
x"00",	-- Hex Addr	6D8D	28045
x"00",	-- Hex Addr	6D8E	28046
x"00",	-- Hex Addr	6D8F	28047
x"00",	-- Hex Addr	6D90	28048
x"00",	-- Hex Addr	6D91	28049
x"00",	-- Hex Addr	6D92	28050
x"00",	-- Hex Addr	6D93	28051
x"00",	-- Hex Addr	6D94	28052
x"00",	-- Hex Addr	6D95	28053
x"00",	-- Hex Addr	6D96	28054
x"00",	-- Hex Addr	6D97	28055
x"00",	-- Hex Addr	6D98	28056
x"00",	-- Hex Addr	6D99	28057
x"00",	-- Hex Addr	6D9A	28058
x"00",	-- Hex Addr	6D9B	28059
x"00",	-- Hex Addr	6D9C	28060
x"00",	-- Hex Addr	6D9D	28061
x"00",	-- Hex Addr	6D9E	28062
x"00",	-- Hex Addr	6D9F	28063
x"00",	-- Hex Addr	6DA0	28064
x"00",	-- Hex Addr	6DA1	28065
x"00",	-- Hex Addr	6DA2	28066
x"00",	-- Hex Addr	6DA3	28067
x"00",	-- Hex Addr	6DA4	28068
x"00",	-- Hex Addr	6DA5	28069
x"00",	-- Hex Addr	6DA6	28070
x"00",	-- Hex Addr	6DA7	28071
x"00",	-- Hex Addr	6DA8	28072
x"00",	-- Hex Addr	6DA9	28073
x"00",	-- Hex Addr	6DAA	28074
x"00",	-- Hex Addr	6DAB	28075
x"00",	-- Hex Addr	6DAC	28076
x"00",	-- Hex Addr	6DAD	28077
x"00",	-- Hex Addr	6DAE	28078
x"00",	-- Hex Addr	6DAF	28079
x"00",	-- Hex Addr	6DB0	28080
x"00",	-- Hex Addr	6DB1	28081
x"00",	-- Hex Addr	6DB2	28082
x"00",	-- Hex Addr	6DB3	28083
x"00",	-- Hex Addr	6DB4	28084
x"00",	-- Hex Addr	6DB5	28085
x"00",	-- Hex Addr	6DB6	28086
x"00",	-- Hex Addr	6DB7	28087
x"00",	-- Hex Addr	6DB8	28088
x"00",	-- Hex Addr	6DB9	28089
x"00",	-- Hex Addr	6DBA	28090
x"00",	-- Hex Addr	6DBB	28091
x"00",	-- Hex Addr	6DBC	28092
x"00",	-- Hex Addr	6DBD	28093
x"00",	-- Hex Addr	6DBE	28094
x"00",	-- Hex Addr	6DBF	28095
x"00",	-- Hex Addr	6DC0	28096
x"00",	-- Hex Addr	6DC1	28097
x"00",	-- Hex Addr	6DC2	28098
x"00",	-- Hex Addr	6DC3	28099
x"00",	-- Hex Addr	6DC4	28100
x"00",	-- Hex Addr	6DC5	28101
x"00",	-- Hex Addr	6DC6	28102
x"00",	-- Hex Addr	6DC7	28103
x"00",	-- Hex Addr	6DC8	28104
x"00",	-- Hex Addr	6DC9	28105
x"00",	-- Hex Addr	6DCA	28106
x"00",	-- Hex Addr	6DCB	28107
x"00",	-- Hex Addr	6DCC	28108
x"00",	-- Hex Addr	6DCD	28109
x"00",	-- Hex Addr	6DCE	28110
x"00",	-- Hex Addr	6DCF	28111
x"00",	-- Hex Addr	6DD0	28112
x"00",	-- Hex Addr	6DD1	28113
x"00",	-- Hex Addr	6DD2	28114
x"00",	-- Hex Addr	6DD3	28115
x"00",	-- Hex Addr	6DD4	28116
x"00",	-- Hex Addr	6DD5	28117
x"00",	-- Hex Addr	6DD6	28118
x"00",	-- Hex Addr	6DD7	28119
x"00",	-- Hex Addr	6DD8	28120
x"00",	-- Hex Addr	6DD9	28121
x"00",	-- Hex Addr	6DDA	28122
x"00",	-- Hex Addr	6DDB	28123
x"00",	-- Hex Addr	6DDC	28124
x"00",	-- Hex Addr	6DDD	28125
x"00",	-- Hex Addr	6DDE	28126
x"00",	-- Hex Addr	6DDF	28127
x"00",	-- Hex Addr	6DE0	28128
x"00",	-- Hex Addr	6DE1	28129
x"00",	-- Hex Addr	6DE2	28130
x"00",	-- Hex Addr	6DE3	28131
x"00",	-- Hex Addr	6DE4	28132
x"00",	-- Hex Addr	6DE5	28133
x"00",	-- Hex Addr	6DE6	28134
x"00",	-- Hex Addr	6DE7	28135
x"00",	-- Hex Addr	6DE8	28136
x"00",	-- Hex Addr	6DE9	28137
x"00",	-- Hex Addr	6DEA	28138
x"00",	-- Hex Addr	6DEB	28139
x"00",	-- Hex Addr	6DEC	28140
x"00",	-- Hex Addr	6DED	28141
x"00",	-- Hex Addr	6DEE	28142
x"00",	-- Hex Addr	6DEF	28143
x"00",	-- Hex Addr	6DF0	28144
x"00",	-- Hex Addr	6DF1	28145
x"00",	-- Hex Addr	6DF2	28146
x"00",	-- Hex Addr	6DF3	28147
x"00",	-- Hex Addr	6DF4	28148
x"00",	-- Hex Addr	6DF5	28149
x"00",	-- Hex Addr	6DF6	28150
x"00",	-- Hex Addr	6DF7	28151
x"00",	-- Hex Addr	6DF8	28152
x"00",	-- Hex Addr	6DF9	28153
x"00",	-- Hex Addr	6DFA	28154
x"00",	-- Hex Addr	6DFB	28155
x"00",	-- Hex Addr	6DFC	28156
x"00",	-- Hex Addr	6DFD	28157
x"00",	-- Hex Addr	6DFE	28158
x"00",	-- Hex Addr	6DFF	28159
x"00",	-- Hex Addr	6E00	28160
x"00",	-- Hex Addr	6E01	28161
x"00",	-- Hex Addr	6E02	28162
x"00",	-- Hex Addr	6E03	28163
x"00",	-- Hex Addr	6E04	28164
x"00",	-- Hex Addr	6E05	28165
x"00",	-- Hex Addr	6E06	28166
x"00",	-- Hex Addr	6E07	28167
x"00",	-- Hex Addr	6E08	28168
x"00",	-- Hex Addr	6E09	28169
x"00",	-- Hex Addr	6E0A	28170
x"00",	-- Hex Addr	6E0B	28171
x"00",	-- Hex Addr	6E0C	28172
x"00",	-- Hex Addr	6E0D	28173
x"00",	-- Hex Addr	6E0E	28174
x"00",	-- Hex Addr	6E0F	28175
x"00",	-- Hex Addr	6E10	28176
x"00",	-- Hex Addr	6E11	28177
x"00",	-- Hex Addr	6E12	28178
x"00",	-- Hex Addr	6E13	28179
x"00",	-- Hex Addr	6E14	28180
x"00",	-- Hex Addr	6E15	28181
x"00",	-- Hex Addr	6E16	28182
x"00",	-- Hex Addr	6E17	28183
x"00",	-- Hex Addr	6E18	28184
x"00",	-- Hex Addr	6E19	28185
x"00",	-- Hex Addr	6E1A	28186
x"00",	-- Hex Addr	6E1B	28187
x"00",	-- Hex Addr	6E1C	28188
x"00",	-- Hex Addr	6E1D	28189
x"00",	-- Hex Addr	6E1E	28190
x"00",	-- Hex Addr	6E1F	28191
x"00",	-- Hex Addr	6E20	28192
x"00",	-- Hex Addr	6E21	28193
x"00",	-- Hex Addr	6E22	28194
x"00",	-- Hex Addr	6E23	28195
x"00",	-- Hex Addr	6E24	28196
x"00",	-- Hex Addr	6E25	28197
x"00",	-- Hex Addr	6E26	28198
x"00",	-- Hex Addr	6E27	28199
x"00",	-- Hex Addr	6E28	28200
x"00",	-- Hex Addr	6E29	28201
x"00",	-- Hex Addr	6E2A	28202
x"00",	-- Hex Addr	6E2B	28203
x"00",	-- Hex Addr	6E2C	28204
x"00",	-- Hex Addr	6E2D	28205
x"00",	-- Hex Addr	6E2E	28206
x"00",	-- Hex Addr	6E2F	28207
x"00",	-- Hex Addr	6E30	28208
x"00",	-- Hex Addr	6E31	28209
x"00",	-- Hex Addr	6E32	28210
x"00",	-- Hex Addr	6E33	28211
x"00",	-- Hex Addr	6E34	28212
x"00",	-- Hex Addr	6E35	28213
x"00",	-- Hex Addr	6E36	28214
x"00",	-- Hex Addr	6E37	28215
x"00",	-- Hex Addr	6E38	28216
x"00",	-- Hex Addr	6E39	28217
x"00",	-- Hex Addr	6E3A	28218
x"00",	-- Hex Addr	6E3B	28219
x"00",	-- Hex Addr	6E3C	28220
x"00",	-- Hex Addr	6E3D	28221
x"00",	-- Hex Addr	6E3E	28222
x"00",	-- Hex Addr	6E3F	28223
x"00",	-- Hex Addr	6E40	28224
x"00",	-- Hex Addr	6E41	28225
x"00",	-- Hex Addr	6E42	28226
x"00",	-- Hex Addr	6E43	28227
x"00",	-- Hex Addr	6E44	28228
x"00",	-- Hex Addr	6E45	28229
x"00",	-- Hex Addr	6E46	28230
x"00",	-- Hex Addr	6E47	28231
x"00",	-- Hex Addr	6E48	28232
x"00",	-- Hex Addr	6E49	28233
x"00",	-- Hex Addr	6E4A	28234
x"00",	-- Hex Addr	6E4B	28235
x"00",	-- Hex Addr	6E4C	28236
x"00",	-- Hex Addr	6E4D	28237
x"00",	-- Hex Addr	6E4E	28238
x"00",	-- Hex Addr	6E4F	28239
x"00",	-- Hex Addr	6E50	28240
x"00",	-- Hex Addr	6E51	28241
x"00",	-- Hex Addr	6E52	28242
x"00",	-- Hex Addr	6E53	28243
x"00",	-- Hex Addr	6E54	28244
x"00",	-- Hex Addr	6E55	28245
x"00",	-- Hex Addr	6E56	28246
x"00",	-- Hex Addr	6E57	28247
x"00",	-- Hex Addr	6E58	28248
x"00",	-- Hex Addr	6E59	28249
x"00",	-- Hex Addr	6E5A	28250
x"00",	-- Hex Addr	6E5B	28251
x"00",	-- Hex Addr	6E5C	28252
x"00",	-- Hex Addr	6E5D	28253
x"00",	-- Hex Addr	6E5E	28254
x"00",	-- Hex Addr	6E5F	28255
x"00",	-- Hex Addr	6E60	28256
x"00",	-- Hex Addr	6E61	28257
x"00",	-- Hex Addr	6E62	28258
x"00",	-- Hex Addr	6E63	28259
x"00",	-- Hex Addr	6E64	28260
x"00",	-- Hex Addr	6E65	28261
x"00",	-- Hex Addr	6E66	28262
x"00",	-- Hex Addr	6E67	28263
x"00",	-- Hex Addr	6E68	28264
x"00",	-- Hex Addr	6E69	28265
x"00",	-- Hex Addr	6E6A	28266
x"00",	-- Hex Addr	6E6B	28267
x"00",	-- Hex Addr	6E6C	28268
x"00",	-- Hex Addr	6E6D	28269
x"00",	-- Hex Addr	6E6E	28270
x"00",	-- Hex Addr	6E6F	28271
x"00",	-- Hex Addr	6E70	28272
x"00",	-- Hex Addr	6E71	28273
x"00",	-- Hex Addr	6E72	28274
x"00",	-- Hex Addr	6E73	28275
x"00",	-- Hex Addr	6E74	28276
x"00",	-- Hex Addr	6E75	28277
x"00",	-- Hex Addr	6E76	28278
x"00",	-- Hex Addr	6E77	28279
x"00",	-- Hex Addr	6E78	28280
x"00",	-- Hex Addr	6E79	28281
x"00",	-- Hex Addr	6E7A	28282
x"00",	-- Hex Addr	6E7B	28283
x"00",	-- Hex Addr	6E7C	28284
x"00",	-- Hex Addr	6E7D	28285
x"00",	-- Hex Addr	6E7E	28286
x"00",	-- Hex Addr	6E7F	28287
x"00",	-- Hex Addr	6E80	28288
x"00",	-- Hex Addr	6E81	28289
x"00",	-- Hex Addr	6E82	28290
x"00",	-- Hex Addr	6E83	28291
x"00",	-- Hex Addr	6E84	28292
x"00",	-- Hex Addr	6E85	28293
x"00",	-- Hex Addr	6E86	28294
x"00",	-- Hex Addr	6E87	28295
x"00",	-- Hex Addr	6E88	28296
x"00",	-- Hex Addr	6E89	28297
x"00",	-- Hex Addr	6E8A	28298
x"00",	-- Hex Addr	6E8B	28299
x"00",	-- Hex Addr	6E8C	28300
x"00",	-- Hex Addr	6E8D	28301
x"00",	-- Hex Addr	6E8E	28302
x"00",	-- Hex Addr	6E8F	28303
x"00",	-- Hex Addr	6E90	28304
x"00",	-- Hex Addr	6E91	28305
x"00",	-- Hex Addr	6E92	28306
x"00",	-- Hex Addr	6E93	28307
x"00",	-- Hex Addr	6E94	28308
x"00",	-- Hex Addr	6E95	28309
x"00",	-- Hex Addr	6E96	28310
x"00",	-- Hex Addr	6E97	28311
x"00",	-- Hex Addr	6E98	28312
x"00",	-- Hex Addr	6E99	28313
x"00",	-- Hex Addr	6E9A	28314
x"00",	-- Hex Addr	6E9B	28315
x"00",	-- Hex Addr	6E9C	28316
x"00",	-- Hex Addr	6E9D	28317
x"00",	-- Hex Addr	6E9E	28318
x"00",	-- Hex Addr	6E9F	28319
x"00",	-- Hex Addr	6EA0	28320
x"00",	-- Hex Addr	6EA1	28321
x"00",	-- Hex Addr	6EA2	28322
x"00",	-- Hex Addr	6EA3	28323
x"00",	-- Hex Addr	6EA4	28324
x"00",	-- Hex Addr	6EA5	28325
x"00",	-- Hex Addr	6EA6	28326
x"00",	-- Hex Addr	6EA7	28327
x"00",	-- Hex Addr	6EA8	28328
x"00",	-- Hex Addr	6EA9	28329
x"00",	-- Hex Addr	6EAA	28330
x"00",	-- Hex Addr	6EAB	28331
x"00",	-- Hex Addr	6EAC	28332
x"00",	-- Hex Addr	6EAD	28333
x"00",	-- Hex Addr	6EAE	28334
x"00",	-- Hex Addr	6EAF	28335
x"00",	-- Hex Addr	6EB0	28336
x"00",	-- Hex Addr	6EB1	28337
x"00",	-- Hex Addr	6EB2	28338
x"00",	-- Hex Addr	6EB3	28339
x"00",	-- Hex Addr	6EB4	28340
x"00",	-- Hex Addr	6EB5	28341
x"00",	-- Hex Addr	6EB6	28342
x"00",	-- Hex Addr	6EB7	28343
x"00",	-- Hex Addr	6EB8	28344
x"00",	-- Hex Addr	6EB9	28345
x"00",	-- Hex Addr	6EBA	28346
x"00",	-- Hex Addr	6EBB	28347
x"00",	-- Hex Addr	6EBC	28348
x"00",	-- Hex Addr	6EBD	28349
x"00",	-- Hex Addr	6EBE	28350
x"00",	-- Hex Addr	6EBF	28351
x"00",	-- Hex Addr	6EC0	28352
x"00",	-- Hex Addr	6EC1	28353
x"00",	-- Hex Addr	6EC2	28354
x"00",	-- Hex Addr	6EC3	28355
x"00",	-- Hex Addr	6EC4	28356
x"00",	-- Hex Addr	6EC5	28357
x"00",	-- Hex Addr	6EC6	28358
x"00",	-- Hex Addr	6EC7	28359
x"00",	-- Hex Addr	6EC8	28360
x"00",	-- Hex Addr	6EC9	28361
x"00",	-- Hex Addr	6ECA	28362
x"00",	-- Hex Addr	6ECB	28363
x"00",	-- Hex Addr	6ECC	28364
x"00",	-- Hex Addr	6ECD	28365
x"00",	-- Hex Addr	6ECE	28366
x"00",	-- Hex Addr	6ECF	28367
x"00",	-- Hex Addr	6ED0	28368
x"00",	-- Hex Addr	6ED1	28369
x"00",	-- Hex Addr	6ED2	28370
x"00",	-- Hex Addr	6ED3	28371
x"00",	-- Hex Addr	6ED4	28372
x"00",	-- Hex Addr	6ED5	28373
x"00",	-- Hex Addr	6ED6	28374
x"00",	-- Hex Addr	6ED7	28375
x"00",	-- Hex Addr	6ED8	28376
x"00",	-- Hex Addr	6ED9	28377
x"00",	-- Hex Addr	6EDA	28378
x"00",	-- Hex Addr	6EDB	28379
x"00",	-- Hex Addr	6EDC	28380
x"00",	-- Hex Addr	6EDD	28381
x"00",	-- Hex Addr	6EDE	28382
x"00",	-- Hex Addr	6EDF	28383
x"00",	-- Hex Addr	6EE0	28384
x"00",	-- Hex Addr	6EE1	28385
x"00",	-- Hex Addr	6EE2	28386
x"00",	-- Hex Addr	6EE3	28387
x"00",	-- Hex Addr	6EE4	28388
x"00",	-- Hex Addr	6EE5	28389
x"00",	-- Hex Addr	6EE6	28390
x"00",	-- Hex Addr	6EE7	28391
x"00",	-- Hex Addr	6EE8	28392
x"00",	-- Hex Addr	6EE9	28393
x"00",	-- Hex Addr	6EEA	28394
x"00",	-- Hex Addr	6EEB	28395
x"00",	-- Hex Addr	6EEC	28396
x"00",	-- Hex Addr	6EED	28397
x"00",	-- Hex Addr	6EEE	28398
x"00",	-- Hex Addr	6EEF	28399
x"00",	-- Hex Addr	6EF0	28400
x"00",	-- Hex Addr	6EF1	28401
x"00",	-- Hex Addr	6EF2	28402
x"00",	-- Hex Addr	6EF3	28403
x"00",	-- Hex Addr	6EF4	28404
x"00",	-- Hex Addr	6EF5	28405
x"00",	-- Hex Addr	6EF6	28406
x"00",	-- Hex Addr	6EF7	28407
x"00",	-- Hex Addr	6EF8	28408
x"00",	-- Hex Addr	6EF9	28409
x"00",	-- Hex Addr	6EFA	28410
x"00",	-- Hex Addr	6EFB	28411
x"00",	-- Hex Addr	6EFC	28412
x"00",	-- Hex Addr	6EFD	28413
x"00",	-- Hex Addr	6EFE	28414
x"00",	-- Hex Addr	6EFF	28415
x"00",	-- Hex Addr	6F00	28416
x"00",	-- Hex Addr	6F01	28417
x"00",	-- Hex Addr	6F02	28418
x"00",	-- Hex Addr	6F03	28419
x"00",	-- Hex Addr	6F04	28420
x"00",	-- Hex Addr	6F05	28421
x"00",	-- Hex Addr	6F06	28422
x"00",	-- Hex Addr	6F07	28423
x"00",	-- Hex Addr	6F08	28424
x"00",	-- Hex Addr	6F09	28425
x"00",	-- Hex Addr	6F0A	28426
x"00",	-- Hex Addr	6F0B	28427
x"00",	-- Hex Addr	6F0C	28428
x"00",	-- Hex Addr	6F0D	28429
x"00",	-- Hex Addr	6F0E	28430
x"00",	-- Hex Addr	6F0F	28431
x"00",	-- Hex Addr	6F10	28432
x"00",	-- Hex Addr	6F11	28433
x"00",	-- Hex Addr	6F12	28434
x"00",	-- Hex Addr	6F13	28435
x"00",	-- Hex Addr	6F14	28436
x"00",	-- Hex Addr	6F15	28437
x"00",	-- Hex Addr	6F16	28438
x"00",	-- Hex Addr	6F17	28439
x"00",	-- Hex Addr	6F18	28440
x"00",	-- Hex Addr	6F19	28441
x"00",	-- Hex Addr	6F1A	28442
x"00",	-- Hex Addr	6F1B	28443
x"00",	-- Hex Addr	6F1C	28444
x"00",	-- Hex Addr	6F1D	28445
x"00",	-- Hex Addr	6F1E	28446
x"00",	-- Hex Addr	6F1F	28447
x"00",	-- Hex Addr	6F20	28448
x"00",	-- Hex Addr	6F21	28449
x"00",	-- Hex Addr	6F22	28450
x"00",	-- Hex Addr	6F23	28451
x"00",	-- Hex Addr	6F24	28452
x"00",	-- Hex Addr	6F25	28453
x"00",	-- Hex Addr	6F26	28454
x"00",	-- Hex Addr	6F27	28455
x"00",	-- Hex Addr	6F28	28456
x"00",	-- Hex Addr	6F29	28457
x"00",	-- Hex Addr	6F2A	28458
x"00",	-- Hex Addr	6F2B	28459
x"00",	-- Hex Addr	6F2C	28460
x"00",	-- Hex Addr	6F2D	28461
x"00",	-- Hex Addr	6F2E	28462
x"00",	-- Hex Addr	6F2F	28463
x"00",	-- Hex Addr	6F30	28464
x"00",	-- Hex Addr	6F31	28465
x"00",	-- Hex Addr	6F32	28466
x"00",	-- Hex Addr	6F33	28467
x"00",	-- Hex Addr	6F34	28468
x"00",	-- Hex Addr	6F35	28469
x"00",	-- Hex Addr	6F36	28470
x"00",	-- Hex Addr	6F37	28471
x"00",	-- Hex Addr	6F38	28472
x"00",	-- Hex Addr	6F39	28473
x"00",	-- Hex Addr	6F3A	28474
x"00",	-- Hex Addr	6F3B	28475
x"00",	-- Hex Addr	6F3C	28476
x"00",	-- Hex Addr	6F3D	28477
x"00",	-- Hex Addr	6F3E	28478
x"00",	-- Hex Addr	6F3F	28479
x"00",	-- Hex Addr	6F40	28480
x"00",	-- Hex Addr	6F41	28481
x"00",	-- Hex Addr	6F42	28482
x"00",	-- Hex Addr	6F43	28483
x"00",	-- Hex Addr	6F44	28484
x"00",	-- Hex Addr	6F45	28485
x"00",	-- Hex Addr	6F46	28486
x"00",	-- Hex Addr	6F47	28487
x"00",	-- Hex Addr	6F48	28488
x"00",	-- Hex Addr	6F49	28489
x"00",	-- Hex Addr	6F4A	28490
x"00",	-- Hex Addr	6F4B	28491
x"00",	-- Hex Addr	6F4C	28492
x"00",	-- Hex Addr	6F4D	28493
x"00",	-- Hex Addr	6F4E	28494
x"00",	-- Hex Addr	6F4F	28495
x"00",	-- Hex Addr	6F50	28496
x"00",	-- Hex Addr	6F51	28497
x"00",	-- Hex Addr	6F52	28498
x"00",	-- Hex Addr	6F53	28499
x"00",	-- Hex Addr	6F54	28500
x"00",	-- Hex Addr	6F55	28501
x"00",	-- Hex Addr	6F56	28502
x"00",	-- Hex Addr	6F57	28503
x"00",	-- Hex Addr	6F58	28504
x"00",	-- Hex Addr	6F59	28505
x"00",	-- Hex Addr	6F5A	28506
x"00",	-- Hex Addr	6F5B	28507
x"00",	-- Hex Addr	6F5C	28508
x"00",	-- Hex Addr	6F5D	28509
x"00",	-- Hex Addr	6F5E	28510
x"00",	-- Hex Addr	6F5F	28511
x"00",	-- Hex Addr	6F60	28512
x"00",	-- Hex Addr	6F61	28513
x"00",	-- Hex Addr	6F62	28514
x"00",	-- Hex Addr	6F63	28515
x"00",	-- Hex Addr	6F64	28516
x"00",	-- Hex Addr	6F65	28517
x"00",	-- Hex Addr	6F66	28518
x"00",	-- Hex Addr	6F67	28519
x"00",	-- Hex Addr	6F68	28520
x"00",	-- Hex Addr	6F69	28521
x"00",	-- Hex Addr	6F6A	28522
x"00",	-- Hex Addr	6F6B	28523
x"00",	-- Hex Addr	6F6C	28524
x"00",	-- Hex Addr	6F6D	28525
x"00",	-- Hex Addr	6F6E	28526
x"00",	-- Hex Addr	6F6F	28527
x"00",	-- Hex Addr	6F70	28528
x"00",	-- Hex Addr	6F71	28529
x"00",	-- Hex Addr	6F72	28530
x"00",	-- Hex Addr	6F73	28531
x"00",	-- Hex Addr	6F74	28532
x"00",	-- Hex Addr	6F75	28533
x"00",	-- Hex Addr	6F76	28534
x"00",	-- Hex Addr	6F77	28535
x"00",	-- Hex Addr	6F78	28536
x"00",	-- Hex Addr	6F79	28537
x"00",	-- Hex Addr	6F7A	28538
x"00",	-- Hex Addr	6F7B	28539
x"00",	-- Hex Addr	6F7C	28540
x"00",	-- Hex Addr	6F7D	28541
x"00",	-- Hex Addr	6F7E	28542
x"00",	-- Hex Addr	6F7F	28543
x"00",	-- Hex Addr	6F80	28544
x"00",	-- Hex Addr	6F81	28545
x"00",	-- Hex Addr	6F82	28546
x"00",	-- Hex Addr	6F83	28547
x"00",	-- Hex Addr	6F84	28548
x"00",	-- Hex Addr	6F85	28549
x"00",	-- Hex Addr	6F86	28550
x"00",	-- Hex Addr	6F87	28551
x"00",	-- Hex Addr	6F88	28552
x"00",	-- Hex Addr	6F89	28553
x"00",	-- Hex Addr	6F8A	28554
x"00",	-- Hex Addr	6F8B	28555
x"00",	-- Hex Addr	6F8C	28556
x"00",	-- Hex Addr	6F8D	28557
x"00",	-- Hex Addr	6F8E	28558
x"00",	-- Hex Addr	6F8F	28559
x"00",	-- Hex Addr	6F90	28560
x"00",	-- Hex Addr	6F91	28561
x"00",	-- Hex Addr	6F92	28562
x"00",	-- Hex Addr	6F93	28563
x"00",	-- Hex Addr	6F94	28564
x"00",	-- Hex Addr	6F95	28565
x"00",	-- Hex Addr	6F96	28566
x"00",	-- Hex Addr	6F97	28567
x"00",	-- Hex Addr	6F98	28568
x"00",	-- Hex Addr	6F99	28569
x"00",	-- Hex Addr	6F9A	28570
x"00",	-- Hex Addr	6F9B	28571
x"00",	-- Hex Addr	6F9C	28572
x"00",	-- Hex Addr	6F9D	28573
x"00",	-- Hex Addr	6F9E	28574
x"00",	-- Hex Addr	6F9F	28575
x"00",	-- Hex Addr	6FA0	28576
x"00",	-- Hex Addr	6FA1	28577
x"00",	-- Hex Addr	6FA2	28578
x"00",	-- Hex Addr	6FA3	28579
x"00",	-- Hex Addr	6FA4	28580
x"00",	-- Hex Addr	6FA5	28581
x"00",	-- Hex Addr	6FA6	28582
x"00",	-- Hex Addr	6FA7	28583
x"00",	-- Hex Addr	6FA8	28584
x"00",	-- Hex Addr	6FA9	28585
x"00",	-- Hex Addr	6FAA	28586
x"00",	-- Hex Addr	6FAB	28587
x"00",	-- Hex Addr	6FAC	28588
x"00",	-- Hex Addr	6FAD	28589
x"00",	-- Hex Addr	6FAE	28590
x"00",	-- Hex Addr	6FAF	28591
x"00",	-- Hex Addr	6FB0	28592
x"00",	-- Hex Addr	6FB1	28593
x"00",	-- Hex Addr	6FB2	28594
x"00",	-- Hex Addr	6FB3	28595
x"00",	-- Hex Addr	6FB4	28596
x"00",	-- Hex Addr	6FB5	28597
x"00",	-- Hex Addr	6FB6	28598
x"00",	-- Hex Addr	6FB7	28599
x"00",	-- Hex Addr	6FB8	28600
x"00",	-- Hex Addr	6FB9	28601
x"00",	-- Hex Addr	6FBA	28602
x"00",	-- Hex Addr	6FBB	28603
x"00",	-- Hex Addr	6FBC	28604
x"00",	-- Hex Addr	6FBD	28605
x"00",	-- Hex Addr	6FBE	28606
x"00",	-- Hex Addr	6FBF	28607
x"00",	-- Hex Addr	6FC0	28608
x"00",	-- Hex Addr	6FC1	28609
x"00",	-- Hex Addr	6FC2	28610
x"00",	-- Hex Addr	6FC3	28611
x"00",	-- Hex Addr	6FC4	28612
x"00",	-- Hex Addr	6FC5	28613
x"00",	-- Hex Addr	6FC6	28614
x"00",	-- Hex Addr	6FC7	28615
x"00",	-- Hex Addr	6FC8	28616
x"00",	-- Hex Addr	6FC9	28617
x"00",	-- Hex Addr	6FCA	28618
x"00",	-- Hex Addr	6FCB	28619
x"00",	-- Hex Addr	6FCC	28620
x"00",	-- Hex Addr	6FCD	28621
x"00",	-- Hex Addr	6FCE	28622
x"00",	-- Hex Addr	6FCF	28623
x"00",	-- Hex Addr	6FD0	28624
x"00",	-- Hex Addr	6FD1	28625
x"00",	-- Hex Addr	6FD2	28626
x"00",	-- Hex Addr	6FD3	28627
x"00",	-- Hex Addr	6FD4	28628
x"00",	-- Hex Addr	6FD5	28629
x"00",	-- Hex Addr	6FD6	28630
x"00",	-- Hex Addr	6FD7	28631
x"00",	-- Hex Addr	6FD8	28632
x"00",	-- Hex Addr	6FD9	28633
x"00",	-- Hex Addr	6FDA	28634
x"00",	-- Hex Addr	6FDB	28635
x"00",	-- Hex Addr	6FDC	28636
x"00",	-- Hex Addr	6FDD	28637
x"00",	-- Hex Addr	6FDE	28638
x"00",	-- Hex Addr	6FDF	28639
x"00",	-- Hex Addr	6FE0	28640
x"00",	-- Hex Addr	6FE1	28641
x"00",	-- Hex Addr	6FE2	28642
x"00",	-- Hex Addr	6FE3	28643
x"00",	-- Hex Addr	6FE4	28644
x"00",	-- Hex Addr	6FE5	28645
x"00",	-- Hex Addr	6FE6	28646
x"00",	-- Hex Addr	6FE7	28647
x"00",	-- Hex Addr	6FE8	28648
x"00",	-- Hex Addr	6FE9	28649
x"00",	-- Hex Addr	6FEA	28650
x"00",	-- Hex Addr	6FEB	28651
x"00",	-- Hex Addr	6FEC	28652
x"00",	-- Hex Addr	6FED	28653
x"00",	-- Hex Addr	6FEE	28654
x"00",	-- Hex Addr	6FEF	28655
x"00",	-- Hex Addr	6FF0	28656
x"00",	-- Hex Addr	6FF1	28657
x"00",	-- Hex Addr	6FF2	28658
x"00",	-- Hex Addr	6FF3	28659
x"00",	-- Hex Addr	6FF4	28660
x"00",	-- Hex Addr	6FF5	28661
x"00",	-- Hex Addr	6FF6	28662
x"00",	-- Hex Addr	6FF7	28663
x"00",	-- Hex Addr	6FF8	28664
x"00",	-- Hex Addr	6FF9	28665
x"00",	-- Hex Addr	6FFA	28666
x"00",	-- Hex Addr	6FFB	28667
x"00",	-- Hex Addr	6FFC	28668
x"00",	-- Hex Addr	6FFD	28669
x"00",	-- Hex Addr	6FFE	28670
x"00",	-- Hex Addr	6FFF	28671
x"00",	-- Hex Addr	7000	28672
x"00",	-- Hex Addr	7001	28673
x"00",	-- Hex Addr	7002	28674
x"00",	-- Hex Addr	7003	28675
x"00",	-- Hex Addr	7004	28676
x"00",	-- Hex Addr	7005	28677
x"00",	-- Hex Addr	7006	28678
x"00",	-- Hex Addr	7007	28679
x"00",	-- Hex Addr	7008	28680
x"00",	-- Hex Addr	7009	28681
x"00",	-- Hex Addr	700A	28682
x"00",	-- Hex Addr	700B	28683
x"00",	-- Hex Addr	700C	28684
x"00",	-- Hex Addr	700D	28685
x"00",	-- Hex Addr	700E	28686
x"00",	-- Hex Addr	700F	28687
x"00",	-- Hex Addr	7010	28688
x"00",	-- Hex Addr	7011	28689
x"00",	-- Hex Addr	7012	28690
x"00",	-- Hex Addr	7013	28691
x"00",	-- Hex Addr	7014	28692
x"00",	-- Hex Addr	7015	28693
x"00",	-- Hex Addr	7016	28694
x"00",	-- Hex Addr	7017	28695
x"00",	-- Hex Addr	7018	28696
x"00",	-- Hex Addr	7019	28697
x"00",	-- Hex Addr	701A	28698
x"00",	-- Hex Addr	701B	28699
x"00",	-- Hex Addr	701C	28700
x"00",	-- Hex Addr	701D	28701
x"00",	-- Hex Addr	701E	28702
x"00",	-- Hex Addr	701F	28703
x"00",	-- Hex Addr	7020	28704
x"00",	-- Hex Addr	7021	28705
x"00",	-- Hex Addr	7022	28706
x"00",	-- Hex Addr	7023	28707
x"00",	-- Hex Addr	7024	28708
x"00",	-- Hex Addr	7025	28709
x"00",	-- Hex Addr	7026	28710
x"00",	-- Hex Addr	7027	28711
x"00",	-- Hex Addr	7028	28712
x"00",	-- Hex Addr	7029	28713
x"00",	-- Hex Addr	702A	28714
x"00",	-- Hex Addr	702B	28715
x"00",	-- Hex Addr	702C	28716
x"00",	-- Hex Addr	702D	28717
x"00",	-- Hex Addr	702E	28718
x"00",	-- Hex Addr	702F	28719
x"00",	-- Hex Addr	7030	28720
x"00",	-- Hex Addr	7031	28721
x"00",	-- Hex Addr	7032	28722
x"00",	-- Hex Addr	7033	28723
x"00",	-- Hex Addr	7034	28724
x"00",	-- Hex Addr	7035	28725
x"00",	-- Hex Addr	7036	28726
x"00",	-- Hex Addr	7037	28727
x"00",	-- Hex Addr	7038	28728
x"00",	-- Hex Addr	7039	28729
x"00",	-- Hex Addr	703A	28730
x"00",	-- Hex Addr	703B	28731
x"00",	-- Hex Addr	703C	28732
x"00",	-- Hex Addr	703D	28733
x"00",	-- Hex Addr	703E	28734
x"00",	-- Hex Addr	703F	28735
x"00",	-- Hex Addr	7040	28736
x"00",	-- Hex Addr	7041	28737
x"00",	-- Hex Addr	7042	28738
x"00",	-- Hex Addr	7043	28739
x"00",	-- Hex Addr	7044	28740
x"00",	-- Hex Addr	7045	28741
x"00",	-- Hex Addr	7046	28742
x"00",	-- Hex Addr	7047	28743
x"00",	-- Hex Addr	7048	28744
x"00",	-- Hex Addr	7049	28745
x"00",	-- Hex Addr	704A	28746
x"00",	-- Hex Addr	704B	28747
x"00",	-- Hex Addr	704C	28748
x"00",	-- Hex Addr	704D	28749
x"00",	-- Hex Addr	704E	28750
x"00",	-- Hex Addr	704F	28751
x"00",	-- Hex Addr	7050	28752
x"00",	-- Hex Addr	7051	28753
x"00",	-- Hex Addr	7052	28754
x"00",	-- Hex Addr	7053	28755
x"00",	-- Hex Addr	7054	28756
x"00",	-- Hex Addr	7055	28757
x"00",	-- Hex Addr	7056	28758
x"00",	-- Hex Addr	7057	28759
x"00",	-- Hex Addr	7058	28760
x"00",	-- Hex Addr	7059	28761
x"00",	-- Hex Addr	705A	28762
x"00",	-- Hex Addr	705B	28763
x"00",	-- Hex Addr	705C	28764
x"00",	-- Hex Addr	705D	28765
x"00",	-- Hex Addr	705E	28766
x"00",	-- Hex Addr	705F	28767
x"00",	-- Hex Addr	7060	28768
x"00",	-- Hex Addr	7061	28769
x"00",	-- Hex Addr	7062	28770
x"00",	-- Hex Addr	7063	28771
x"00",	-- Hex Addr	7064	28772
x"00",	-- Hex Addr	7065	28773
x"00",	-- Hex Addr	7066	28774
x"00",	-- Hex Addr	7067	28775
x"00",	-- Hex Addr	7068	28776
x"00",	-- Hex Addr	7069	28777
x"00",	-- Hex Addr	706A	28778
x"00",	-- Hex Addr	706B	28779
x"00",	-- Hex Addr	706C	28780
x"00",	-- Hex Addr	706D	28781
x"00",	-- Hex Addr	706E	28782
x"00",	-- Hex Addr	706F	28783
x"00",	-- Hex Addr	7070	28784
x"00",	-- Hex Addr	7071	28785
x"00",	-- Hex Addr	7072	28786
x"00",	-- Hex Addr	7073	28787
x"00",	-- Hex Addr	7074	28788
x"00",	-- Hex Addr	7075	28789
x"00",	-- Hex Addr	7076	28790
x"00",	-- Hex Addr	7077	28791
x"00",	-- Hex Addr	7078	28792
x"00",	-- Hex Addr	7079	28793
x"00",	-- Hex Addr	707A	28794
x"00",	-- Hex Addr	707B	28795
x"00",	-- Hex Addr	707C	28796
x"00",	-- Hex Addr	707D	28797
x"00",	-- Hex Addr	707E	28798
x"00",	-- Hex Addr	707F	28799
x"00",	-- Hex Addr	7080	28800
x"00",	-- Hex Addr	7081	28801
x"00",	-- Hex Addr	7082	28802
x"00",	-- Hex Addr	7083	28803
x"00",	-- Hex Addr	7084	28804
x"00",	-- Hex Addr	7085	28805
x"00",	-- Hex Addr	7086	28806
x"00",	-- Hex Addr	7087	28807
x"00",	-- Hex Addr	7088	28808
x"00",	-- Hex Addr	7089	28809
x"00",	-- Hex Addr	708A	28810
x"00",	-- Hex Addr	708B	28811
x"00",	-- Hex Addr	708C	28812
x"00",	-- Hex Addr	708D	28813
x"00",	-- Hex Addr	708E	28814
x"00",	-- Hex Addr	708F	28815
x"00",	-- Hex Addr	7090	28816
x"00",	-- Hex Addr	7091	28817
x"00",	-- Hex Addr	7092	28818
x"00",	-- Hex Addr	7093	28819
x"00",	-- Hex Addr	7094	28820
x"00",	-- Hex Addr	7095	28821
x"00",	-- Hex Addr	7096	28822
x"00",	-- Hex Addr	7097	28823
x"00",	-- Hex Addr	7098	28824
x"00",	-- Hex Addr	7099	28825
x"00",	-- Hex Addr	709A	28826
x"00",	-- Hex Addr	709B	28827
x"00",	-- Hex Addr	709C	28828
x"00",	-- Hex Addr	709D	28829
x"00",	-- Hex Addr	709E	28830
x"00",	-- Hex Addr	709F	28831
x"00",	-- Hex Addr	70A0	28832
x"00",	-- Hex Addr	70A1	28833
x"00",	-- Hex Addr	70A2	28834
x"00",	-- Hex Addr	70A3	28835
x"00",	-- Hex Addr	70A4	28836
x"00",	-- Hex Addr	70A5	28837
x"00",	-- Hex Addr	70A6	28838
x"00",	-- Hex Addr	70A7	28839
x"00",	-- Hex Addr	70A8	28840
x"00",	-- Hex Addr	70A9	28841
x"00",	-- Hex Addr	70AA	28842
x"00",	-- Hex Addr	70AB	28843
x"00",	-- Hex Addr	70AC	28844
x"00",	-- Hex Addr	70AD	28845
x"00",	-- Hex Addr	70AE	28846
x"00",	-- Hex Addr	70AF	28847
x"00",	-- Hex Addr	70B0	28848
x"00",	-- Hex Addr	70B1	28849
x"00",	-- Hex Addr	70B2	28850
x"00",	-- Hex Addr	70B3	28851
x"00",	-- Hex Addr	70B4	28852
x"00",	-- Hex Addr	70B5	28853
x"00",	-- Hex Addr	70B6	28854
x"00",	-- Hex Addr	70B7	28855
x"00",	-- Hex Addr	70B8	28856
x"00",	-- Hex Addr	70B9	28857
x"00",	-- Hex Addr	70BA	28858
x"00",	-- Hex Addr	70BB	28859
x"00",	-- Hex Addr	70BC	28860
x"00",	-- Hex Addr	70BD	28861
x"00",	-- Hex Addr	70BE	28862
x"00",	-- Hex Addr	70BF	28863
x"00",	-- Hex Addr	70C0	28864
x"00",	-- Hex Addr	70C1	28865
x"00",	-- Hex Addr	70C2	28866
x"00",	-- Hex Addr	70C3	28867
x"00",	-- Hex Addr	70C4	28868
x"00",	-- Hex Addr	70C5	28869
x"00",	-- Hex Addr	70C6	28870
x"00",	-- Hex Addr	70C7	28871
x"00",	-- Hex Addr	70C8	28872
x"00",	-- Hex Addr	70C9	28873
x"00",	-- Hex Addr	70CA	28874
x"00",	-- Hex Addr	70CB	28875
x"00",	-- Hex Addr	70CC	28876
x"00",	-- Hex Addr	70CD	28877
x"00",	-- Hex Addr	70CE	28878
x"00",	-- Hex Addr	70CF	28879
x"00",	-- Hex Addr	70D0	28880
x"00",	-- Hex Addr	70D1	28881
x"00",	-- Hex Addr	70D2	28882
x"00",	-- Hex Addr	70D3	28883
x"00",	-- Hex Addr	70D4	28884
x"00",	-- Hex Addr	70D5	28885
x"00",	-- Hex Addr	70D6	28886
x"00",	-- Hex Addr	70D7	28887
x"00",	-- Hex Addr	70D8	28888
x"00",	-- Hex Addr	70D9	28889
x"00",	-- Hex Addr	70DA	28890
x"00",	-- Hex Addr	70DB	28891
x"00",	-- Hex Addr	70DC	28892
x"00",	-- Hex Addr	70DD	28893
x"00",	-- Hex Addr	70DE	28894
x"00",	-- Hex Addr	70DF	28895
x"00",	-- Hex Addr	70E0	28896
x"00",	-- Hex Addr	70E1	28897
x"00",	-- Hex Addr	70E2	28898
x"00",	-- Hex Addr	70E3	28899
x"00",	-- Hex Addr	70E4	28900
x"00",	-- Hex Addr	70E5	28901
x"00",	-- Hex Addr	70E6	28902
x"00",	-- Hex Addr	70E7	28903
x"00",	-- Hex Addr	70E8	28904
x"00",	-- Hex Addr	70E9	28905
x"00",	-- Hex Addr	70EA	28906
x"00",	-- Hex Addr	70EB	28907
x"00",	-- Hex Addr	70EC	28908
x"00",	-- Hex Addr	70ED	28909
x"00",	-- Hex Addr	70EE	28910
x"00",	-- Hex Addr	70EF	28911
x"00",	-- Hex Addr	70F0	28912
x"00",	-- Hex Addr	70F1	28913
x"00",	-- Hex Addr	70F2	28914
x"00",	-- Hex Addr	70F3	28915
x"00",	-- Hex Addr	70F4	28916
x"00",	-- Hex Addr	70F5	28917
x"00",	-- Hex Addr	70F6	28918
x"00",	-- Hex Addr	70F7	28919
x"00",	-- Hex Addr	70F8	28920
x"00",	-- Hex Addr	70F9	28921
x"00",	-- Hex Addr	70FA	28922
x"00",	-- Hex Addr	70FB	28923
x"00",	-- Hex Addr	70FC	28924
x"00",	-- Hex Addr	70FD	28925
x"00",	-- Hex Addr	70FE	28926
x"00",	-- Hex Addr	70FF	28927
x"00",	-- Hex Addr	7100	28928
x"00",	-- Hex Addr	7101	28929
x"00",	-- Hex Addr	7102	28930
x"00",	-- Hex Addr	7103	28931
x"00",	-- Hex Addr	7104	28932
x"00",	-- Hex Addr	7105	28933
x"00",	-- Hex Addr	7106	28934
x"00",	-- Hex Addr	7107	28935
x"00",	-- Hex Addr	7108	28936
x"00",	-- Hex Addr	7109	28937
x"00",	-- Hex Addr	710A	28938
x"00",	-- Hex Addr	710B	28939
x"00",	-- Hex Addr	710C	28940
x"00",	-- Hex Addr	710D	28941
x"00",	-- Hex Addr	710E	28942
x"00",	-- Hex Addr	710F	28943
x"00",	-- Hex Addr	7110	28944
x"00",	-- Hex Addr	7111	28945
x"00",	-- Hex Addr	7112	28946
x"00",	-- Hex Addr	7113	28947
x"00",	-- Hex Addr	7114	28948
x"00",	-- Hex Addr	7115	28949
x"00",	-- Hex Addr	7116	28950
x"00",	-- Hex Addr	7117	28951
x"00",	-- Hex Addr	7118	28952
x"00",	-- Hex Addr	7119	28953
x"00",	-- Hex Addr	711A	28954
x"00",	-- Hex Addr	711B	28955
x"00",	-- Hex Addr	711C	28956
x"00",	-- Hex Addr	711D	28957
x"00",	-- Hex Addr	711E	28958
x"00",	-- Hex Addr	711F	28959
x"00",	-- Hex Addr	7120	28960
x"00",	-- Hex Addr	7121	28961
x"00",	-- Hex Addr	7122	28962
x"00",	-- Hex Addr	7123	28963
x"00",	-- Hex Addr	7124	28964
x"00",	-- Hex Addr	7125	28965
x"00",	-- Hex Addr	7126	28966
x"00",	-- Hex Addr	7127	28967
x"00",	-- Hex Addr	7128	28968
x"00",	-- Hex Addr	7129	28969
x"00",	-- Hex Addr	712A	28970
x"00",	-- Hex Addr	712B	28971
x"00",	-- Hex Addr	712C	28972
x"00",	-- Hex Addr	712D	28973
x"00",	-- Hex Addr	712E	28974
x"00",	-- Hex Addr	712F	28975
x"00",	-- Hex Addr	7130	28976
x"00",	-- Hex Addr	7131	28977
x"00",	-- Hex Addr	7132	28978
x"00",	-- Hex Addr	7133	28979
x"00",	-- Hex Addr	7134	28980
x"00",	-- Hex Addr	7135	28981
x"00",	-- Hex Addr	7136	28982
x"00",	-- Hex Addr	7137	28983
x"00",	-- Hex Addr	7138	28984
x"00",	-- Hex Addr	7139	28985
x"00",	-- Hex Addr	713A	28986
x"00",	-- Hex Addr	713B	28987
x"00",	-- Hex Addr	713C	28988
x"00",	-- Hex Addr	713D	28989
x"00",	-- Hex Addr	713E	28990
x"00",	-- Hex Addr	713F	28991
x"00",	-- Hex Addr	7140	28992
x"00",	-- Hex Addr	7141	28993
x"00",	-- Hex Addr	7142	28994
x"00",	-- Hex Addr	7143	28995
x"00",	-- Hex Addr	7144	28996
x"00",	-- Hex Addr	7145	28997
x"00",	-- Hex Addr	7146	28998
x"00",	-- Hex Addr	7147	28999
x"00",	-- Hex Addr	7148	29000
x"00",	-- Hex Addr	7149	29001
x"00",	-- Hex Addr	714A	29002
x"00",	-- Hex Addr	714B	29003
x"00",	-- Hex Addr	714C	29004
x"00",	-- Hex Addr	714D	29005
x"00",	-- Hex Addr	714E	29006
x"00",	-- Hex Addr	714F	29007
x"00",	-- Hex Addr	7150	29008
x"00",	-- Hex Addr	7151	29009
x"00",	-- Hex Addr	7152	29010
x"00",	-- Hex Addr	7153	29011
x"00",	-- Hex Addr	7154	29012
x"00",	-- Hex Addr	7155	29013
x"00",	-- Hex Addr	7156	29014
x"00",	-- Hex Addr	7157	29015
x"00",	-- Hex Addr	7158	29016
x"00",	-- Hex Addr	7159	29017
x"00",	-- Hex Addr	715A	29018
x"00",	-- Hex Addr	715B	29019
x"00",	-- Hex Addr	715C	29020
x"00",	-- Hex Addr	715D	29021
x"00",	-- Hex Addr	715E	29022
x"00",	-- Hex Addr	715F	29023
x"00",	-- Hex Addr	7160	29024
x"00",	-- Hex Addr	7161	29025
x"00",	-- Hex Addr	7162	29026
x"00",	-- Hex Addr	7163	29027
x"00",	-- Hex Addr	7164	29028
x"00",	-- Hex Addr	7165	29029
x"00",	-- Hex Addr	7166	29030
x"00",	-- Hex Addr	7167	29031
x"00",	-- Hex Addr	7168	29032
x"00",	-- Hex Addr	7169	29033
x"00",	-- Hex Addr	716A	29034
x"00",	-- Hex Addr	716B	29035
x"00",	-- Hex Addr	716C	29036
x"00",	-- Hex Addr	716D	29037
x"00",	-- Hex Addr	716E	29038
x"00",	-- Hex Addr	716F	29039
x"00",	-- Hex Addr	7170	29040
x"00",	-- Hex Addr	7171	29041
x"00",	-- Hex Addr	7172	29042
x"00",	-- Hex Addr	7173	29043
x"00",	-- Hex Addr	7174	29044
x"00",	-- Hex Addr	7175	29045
x"00",	-- Hex Addr	7176	29046
x"00",	-- Hex Addr	7177	29047
x"00",	-- Hex Addr	7178	29048
x"00",	-- Hex Addr	7179	29049
x"00",	-- Hex Addr	717A	29050
x"00",	-- Hex Addr	717B	29051
x"00",	-- Hex Addr	717C	29052
x"00",	-- Hex Addr	717D	29053
x"00",	-- Hex Addr	717E	29054
x"00",	-- Hex Addr	717F	29055
x"00",	-- Hex Addr	7180	29056
x"00",	-- Hex Addr	7181	29057
x"00",	-- Hex Addr	7182	29058
x"00",	-- Hex Addr	7183	29059
x"00",	-- Hex Addr	7184	29060
x"00",	-- Hex Addr	7185	29061
x"00",	-- Hex Addr	7186	29062
x"00",	-- Hex Addr	7187	29063
x"00",	-- Hex Addr	7188	29064
x"00",	-- Hex Addr	7189	29065
x"00",	-- Hex Addr	718A	29066
x"00",	-- Hex Addr	718B	29067
x"00",	-- Hex Addr	718C	29068
x"00",	-- Hex Addr	718D	29069
x"00",	-- Hex Addr	718E	29070
x"00",	-- Hex Addr	718F	29071
x"00",	-- Hex Addr	7190	29072
x"00",	-- Hex Addr	7191	29073
x"00",	-- Hex Addr	7192	29074
x"00",	-- Hex Addr	7193	29075
x"00",	-- Hex Addr	7194	29076
x"00",	-- Hex Addr	7195	29077
x"00",	-- Hex Addr	7196	29078
x"00",	-- Hex Addr	7197	29079
x"00",	-- Hex Addr	7198	29080
x"00",	-- Hex Addr	7199	29081
x"00",	-- Hex Addr	719A	29082
x"00",	-- Hex Addr	719B	29083
x"00",	-- Hex Addr	719C	29084
x"00",	-- Hex Addr	719D	29085
x"00",	-- Hex Addr	719E	29086
x"00",	-- Hex Addr	719F	29087
x"00",	-- Hex Addr	71A0	29088
x"00",	-- Hex Addr	71A1	29089
x"00",	-- Hex Addr	71A2	29090
x"00",	-- Hex Addr	71A3	29091
x"00",	-- Hex Addr	71A4	29092
x"00",	-- Hex Addr	71A5	29093
x"00",	-- Hex Addr	71A6	29094
x"00",	-- Hex Addr	71A7	29095
x"00",	-- Hex Addr	71A8	29096
x"00",	-- Hex Addr	71A9	29097
x"00",	-- Hex Addr	71AA	29098
x"00",	-- Hex Addr	71AB	29099
x"00",	-- Hex Addr	71AC	29100
x"00",	-- Hex Addr	71AD	29101
x"00",	-- Hex Addr	71AE	29102
x"00",	-- Hex Addr	71AF	29103
x"00",	-- Hex Addr	71B0	29104
x"00",	-- Hex Addr	71B1	29105
x"00",	-- Hex Addr	71B2	29106
x"00",	-- Hex Addr	71B3	29107
x"00",	-- Hex Addr	71B4	29108
x"00",	-- Hex Addr	71B5	29109
x"00",	-- Hex Addr	71B6	29110
x"00",	-- Hex Addr	71B7	29111
x"00",	-- Hex Addr	71B8	29112
x"00",	-- Hex Addr	71B9	29113
x"00",	-- Hex Addr	71BA	29114
x"00",	-- Hex Addr	71BB	29115
x"00",	-- Hex Addr	71BC	29116
x"00",	-- Hex Addr	71BD	29117
x"00",	-- Hex Addr	71BE	29118
x"00",	-- Hex Addr	71BF	29119
x"00",	-- Hex Addr	71C0	29120
x"00",	-- Hex Addr	71C1	29121
x"00",	-- Hex Addr	71C2	29122
x"00",	-- Hex Addr	71C3	29123
x"00",	-- Hex Addr	71C4	29124
x"00",	-- Hex Addr	71C5	29125
x"00",	-- Hex Addr	71C6	29126
x"00",	-- Hex Addr	71C7	29127
x"00",	-- Hex Addr	71C8	29128
x"00",	-- Hex Addr	71C9	29129
x"00",	-- Hex Addr	71CA	29130
x"00",	-- Hex Addr	71CB	29131
x"00",	-- Hex Addr	71CC	29132
x"00",	-- Hex Addr	71CD	29133
x"00",	-- Hex Addr	71CE	29134
x"00",	-- Hex Addr	71CF	29135
x"00",	-- Hex Addr	71D0	29136
x"00",	-- Hex Addr	71D1	29137
x"00",	-- Hex Addr	71D2	29138
x"00",	-- Hex Addr	71D3	29139
x"00",	-- Hex Addr	71D4	29140
x"00",	-- Hex Addr	71D5	29141
x"00",	-- Hex Addr	71D6	29142
x"00",	-- Hex Addr	71D7	29143
x"00",	-- Hex Addr	71D8	29144
x"00",	-- Hex Addr	71D9	29145
x"00",	-- Hex Addr	71DA	29146
x"00",	-- Hex Addr	71DB	29147
x"00",	-- Hex Addr	71DC	29148
x"00",	-- Hex Addr	71DD	29149
x"00",	-- Hex Addr	71DE	29150
x"00",	-- Hex Addr	71DF	29151
x"00",	-- Hex Addr	71E0	29152
x"00",	-- Hex Addr	71E1	29153
x"00",	-- Hex Addr	71E2	29154
x"00",	-- Hex Addr	71E3	29155
x"00",	-- Hex Addr	71E4	29156
x"00",	-- Hex Addr	71E5	29157
x"00",	-- Hex Addr	71E6	29158
x"00",	-- Hex Addr	71E7	29159
x"00",	-- Hex Addr	71E8	29160
x"00",	-- Hex Addr	71E9	29161
x"00",	-- Hex Addr	71EA	29162
x"00",	-- Hex Addr	71EB	29163
x"00",	-- Hex Addr	71EC	29164
x"00",	-- Hex Addr	71ED	29165
x"00",	-- Hex Addr	71EE	29166
x"00",	-- Hex Addr	71EF	29167
x"00",	-- Hex Addr	71F0	29168
x"00",	-- Hex Addr	71F1	29169
x"00",	-- Hex Addr	71F2	29170
x"00",	-- Hex Addr	71F3	29171
x"00",	-- Hex Addr	71F4	29172
x"00",	-- Hex Addr	71F5	29173
x"00",	-- Hex Addr	71F6	29174
x"00",	-- Hex Addr	71F7	29175
x"00",	-- Hex Addr	71F8	29176
x"00",	-- Hex Addr	71F9	29177
x"00",	-- Hex Addr	71FA	29178
x"00",	-- Hex Addr	71FB	29179
x"00",	-- Hex Addr	71FC	29180
x"00",	-- Hex Addr	71FD	29181
x"00",	-- Hex Addr	71FE	29182
x"00",	-- Hex Addr	71FF	29183
x"00",	-- Hex Addr	7200	29184
x"00",	-- Hex Addr	7201	29185
x"00",	-- Hex Addr	7202	29186
x"00",	-- Hex Addr	7203	29187
x"00",	-- Hex Addr	7204	29188
x"00",	-- Hex Addr	7205	29189
x"00",	-- Hex Addr	7206	29190
x"00",	-- Hex Addr	7207	29191
x"00",	-- Hex Addr	7208	29192
x"00",	-- Hex Addr	7209	29193
x"00",	-- Hex Addr	720A	29194
x"00",	-- Hex Addr	720B	29195
x"00",	-- Hex Addr	720C	29196
x"00",	-- Hex Addr	720D	29197
x"00",	-- Hex Addr	720E	29198
x"00",	-- Hex Addr	720F	29199
x"00",	-- Hex Addr	7210	29200
x"00",	-- Hex Addr	7211	29201
x"00",	-- Hex Addr	7212	29202
x"00",	-- Hex Addr	7213	29203
x"00",	-- Hex Addr	7214	29204
x"00",	-- Hex Addr	7215	29205
x"00",	-- Hex Addr	7216	29206
x"00",	-- Hex Addr	7217	29207
x"00",	-- Hex Addr	7218	29208
x"00",	-- Hex Addr	7219	29209
x"00",	-- Hex Addr	721A	29210
x"00",	-- Hex Addr	721B	29211
x"00",	-- Hex Addr	721C	29212
x"00",	-- Hex Addr	721D	29213
x"00",	-- Hex Addr	721E	29214
x"00",	-- Hex Addr	721F	29215
x"00",	-- Hex Addr	7220	29216
x"00",	-- Hex Addr	7221	29217
x"00",	-- Hex Addr	7222	29218
x"00",	-- Hex Addr	7223	29219
x"00",	-- Hex Addr	7224	29220
x"00",	-- Hex Addr	7225	29221
x"00",	-- Hex Addr	7226	29222
x"00",	-- Hex Addr	7227	29223
x"00",	-- Hex Addr	7228	29224
x"00",	-- Hex Addr	7229	29225
x"00",	-- Hex Addr	722A	29226
x"00",	-- Hex Addr	722B	29227
x"00",	-- Hex Addr	722C	29228
x"00",	-- Hex Addr	722D	29229
x"00",	-- Hex Addr	722E	29230
x"00",	-- Hex Addr	722F	29231
x"00",	-- Hex Addr	7230	29232
x"00",	-- Hex Addr	7231	29233
x"00",	-- Hex Addr	7232	29234
x"00",	-- Hex Addr	7233	29235
x"00",	-- Hex Addr	7234	29236
x"00",	-- Hex Addr	7235	29237
x"00",	-- Hex Addr	7236	29238
x"00",	-- Hex Addr	7237	29239
x"00",	-- Hex Addr	7238	29240
x"00",	-- Hex Addr	7239	29241
x"00",	-- Hex Addr	723A	29242
x"00",	-- Hex Addr	723B	29243
x"00",	-- Hex Addr	723C	29244
x"00",	-- Hex Addr	723D	29245
x"00",	-- Hex Addr	723E	29246
x"00",	-- Hex Addr	723F	29247
x"00",	-- Hex Addr	7240	29248
x"00",	-- Hex Addr	7241	29249
x"00",	-- Hex Addr	7242	29250
x"00",	-- Hex Addr	7243	29251
x"00",	-- Hex Addr	7244	29252
x"00",	-- Hex Addr	7245	29253
x"00",	-- Hex Addr	7246	29254
x"00",	-- Hex Addr	7247	29255
x"00",	-- Hex Addr	7248	29256
x"00",	-- Hex Addr	7249	29257
x"00",	-- Hex Addr	724A	29258
x"00",	-- Hex Addr	724B	29259
x"00",	-- Hex Addr	724C	29260
x"00",	-- Hex Addr	724D	29261
x"00",	-- Hex Addr	724E	29262
x"00",	-- Hex Addr	724F	29263
x"00",	-- Hex Addr	7250	29264
x"00",	-- Hex Addr	7251	29265
x"00",	-- Hex Addr	7252	29266
x"00",	-- Hex Addr	7253	29267
x"00",	-- Hex Addr	7254	29268
x"00",	-- Hex Addr	7255	29269
x"00",	-- Hex Addr	7256	29270
x"00",	-- Hex Addr	7257	29271
x"00",	-- Hex Addr	7258	29272
x"00",	-- Hex Addr	7259	29273
x"00",	-- Hex Addr	725A	29274
x"00",	-- Hex Addr	725B	29275
x"00",	-- Hex Addr	725C	29276
x"00",	-- Hex Addr	725D	29277
x"00",	-- Hex Addr	725E	29278
x"00",	-- Hex Addr	725F	29279
x"00",	-- Hex Addr	7260	29280
x"00",	-- Hex Addr	7261	29281
x"00",	-- Hex Addr	7262	29282
x"00",	-- Hex Addr	7263	29283
x"00",	-- Hex Addr	7264	29284
x"00",	-- Hex Addr	7265	29285
x"00",	-- Hex Addr	7266	29286
x"00",	-- Hex Addr	7267	29287
x"00",	-- Hex Addr	7268	29288
x"00",	-- Hex Addr	7269	29289
x"00",	-- Hex Addr	726A	29290
x"00",	-- Hex Addr	726B	29291
x"00",	-- Hex Addr	726C	29292
x"00",	-- Hex Addr	726D	29293
x"00",	-- Hex Addr	726E	29294
x"00",	-- Hex Addr	726F	29295
x"00",	-- Hex Addr	7270	29296
x"00",	-- Hex Addr	7271	29297
x"00",	-- Hex Addr	7272	29298
x"00",	-- Hex Addr	7273	29299
x"00",	-- Hex Addr	7274	29300
x"00",	-- Hex Addr	7275	29301
x"00",	-- Hex Addr	7276	29302
x"00",	-- Hex Addr	7277	29303
x"00",	-- Hex Addr	7278	29304
x"00",	-- Hex Addr	7279	29305
x"00",	-- Hex Addr	727A	29306
x"00",	-- Hex Addr	727B	29307
x"00",	-- Hex Addr	727C	29308
x"00",	-- Hex Addr	727D	29309
x"00",	-- Hex Addr	727E	29310
x"00",	-- Hex Addr	727F	29311
x"00",	-- Hex Addr	7280	29312
x"00",	-- Hex Addr	7281	29313
x"00",	-- Hex Addr	7282	29314
x"00",	-- Hex Addr	7283	29315
x"00",	-- Hex Addr	7284	29316
x"00",	-- Hex Addr	7285	29317
x"00",	-- Hex Addr	7286	29318
x"00",	-- Hex Addr	7287	29319
x"00",	-- Hex Addr	7288	29320
x"00",	-- Hex Addr	7289	29321
x"00",	-- Hex Addr	728A	29322
x"00",	-- Hex Addr	728B	29323
x"00",	-- Hex Addr	728C	29324
x"00",	-- Hex Addr	728D	29325
x"00",	-- Hex Addr	728E	29326
x"00",	-- Hex Addr	728F	29327
x"00",	-- Hex Addr	7290	29328
x"00",	-- Hex Addr	7291	29329
x"00",	-- Hex Addr	7292	29330
x"00",	-- Hex Addr	7293	29331
x"00",	-- Hex Addr	7294	29332
x"00",	-- Hex Addr	7295	29333
x"00",	-- Hex Addr	7296	29334
x"00",	-- Hex Addr	7297	29335
x"00",	-- Hex Addr	7298	29336
x"00",	-- Hex Addr	7299	29337
x"00",	-- Hex Addr	729A	29338
x"00",	-- Hex Addr	729B	29339
x"00",	-- Hex Addr	729C	29340
x"00",	-- Hex Addr	729D	29341
x"00",	-- Hex Addr	729E	29342
x"00",	-- Hex Addr	729F	29343
x"00",	-- Hex Addr	72A0	29344
x"00",	-- Hex Addr	72A1	29345
x"00",	-- Hex Addr	72A2	29346
x"00",	-- Hex Addr	72A3	29347
x"00",	-- Hex Addr	72A4	29348
x"00",	-- Hex Addr	72A5	29349
x"00",	-- Hex Addr	72A6	29350
x"00",	-- Hex Addr	72A7	29351
x"00",	-- Hex Addr	72A8	29352
x"00",	-- Hex Addr	72A9	29353
x"00",	-- Hex Addr	72AA	29354
x"00",	-- Hex Addr	72AB	29355
x"00",	-- Hex Addr	72AC	29356
x"00",	-- Hex Addr	72AD	29357
x"00",	-- Hex Addr	72AE	29358
x"00",	-- Hex Addr	72AF	29359
x"00",	-- Hex Addr	72B0	29360
x"00",	-- Hex Addr	72B1	29361
x"00",	-- Hex Addr	72B2	29362
x"00",	-- Hex Addr	72B3	29363
x"00",	-- Hex Addr	72B4	29364
x"00",	-- Hex Addr	72B5	29365
x"00",	-- Hex Addr	72B6	29366
x"00",	-- Hex Addr	72B7	29367
x"00",	-- Hex Addr	72B8	29368
x"00",	-- Hex Addr	72B9	29369
x"00",	-- Hex Addr	72BA	29370
x"00",	-- Hex Addr	72BB	29371
x"00",	-- Hex Addr	72BC	29372
x"00",	-- Hex Addr	72BD	29373
x"00",	-- Hex Addr	72BE	29374
x"00",	-- Hex Addr	72BF	29375
x"00",	-- Hex Addr	72C0	29376
x"00",	-- Hex Addr	72C1	29377
x"00",	-- Hex Addr	72C2	29378
x"00",	-- Hex Addr	72C3	29379
x"00",	-- Hex Addr	72C4	29380
x"00",	-- Hex Addr	72C5	29381
x"00",	-- Hex Addr	72C6	29382
x"00",	-- Hex Addr	72C7	29383
x"00",	-- Hex Addr	72C8	29384
x"00",	-- Hex Addr	72C9	29385
x"00",	-- Hex Addr	72CA	29386
x"00",	-- Hex Addr	72CB	29387
x"00",	-- Hex Addr	72CC	29388
x"00",	-- Hex Addr	72CD	29389
x"00",	-- Hex Addr	72CE	29390
x"00",	-- Hex Addr	72CF	29391
x"00",	-- Hex Addr	72D0	29392
x"00",	-- Hex Addr	72D1	29393
x"00",	-- Hex Addr	72D2	29394
x"00",	-- Hex Addr	72D3	29395
x"00",	-- Hex Addr	72D4	29396
x"00",	-- Hex Addr	72D5	29397
x"00",	-- Hex Addr	72D6	29398
x"00",	-- Hex Addr	72D7	29399
x"00",	-- Hex Addr	72D8	29400
x"00",	-- Hex Addr	72D9	29401
x"00",	-- Hex Addr	72DA	29402
x"00",	-- Hex Addr	72DB	29403
x"00",	-- Hex Addr	72DC	29404
x"00",	-- Hex Addr	72DD	29405
x"00",	-- Hex Addr	72DE	29406
x"00",	-- Hex Addr	72DF	29407
x"00",	-- Hex Addr	72E0	29408
x"00",	-- Hex Addr	72E1	29409
x"00",	-- Hex Addr	72E2	29410
x"00",	-- Hex Addr	72E3	29411
x"00",	-- Hex Addr	72E4	29412
x"00",	-- Hex Addr	72E5	29413
x"00",	-- Hex Addr	72E6	29414
x"00",	-- Hex Addr	72E7	29415
x"00",	-- Hex Addr	72E8	29416
x"00",	-- Hex Addr	72E9	29417
x"00",	-- Hex Addr	72EA	29418
x"00",	-- Hex Addr	72EB	29419
x"00",	-- Hex Addr	72EC	29420
x"00",	-- Hex Addr	72ED	29421
x"00",	-- Hex Addr	72EE	29422
x"00",	-- Hex Addr	72EF	29423
x"00",	-- Hex Addr	72F0	29424
x"00",	-- Hex Addr	72F1	29425
x"00",	-- Hex Addr	72F2	29426
x"00",	-- Hex Addr	72F3	29427
x"00",	-- Hex Addr	72F4	29428
x"00",	-- Hex Addr	72F5	29429
x"00",	-- Hex Addr	72F6	29430
x"00",	-- Hex Addr	72F7	29431
x"00",	-- Hex Addr	72F8	29432
x"00",	-- Hex Addr	72F9	29433
x"00",	-- Hex Addr	72FA	29434
x"00",	-- Hex Addr	72FB	29435
x"00",	-- Hex Addr	72FC	29436
x"00",	-- Hex Addr	72FD	29437
x"00",	-- Hex Addr	72FE	29438
x"00",	-- Hex Addr	72FF	29439
x"00",	-- Hex Addr	7300	29440
x"00",	-- Hex Addr	7301	29441
x"00",	-- Hex Addr	7302	29442
x"00",	-- Hex Addr	7303	29443
x"00",	-- Hex Addr	7304	29444
x"00",	-- Hex Addr	7305	29445
x"00",	-- Hex Addr	7306	29446
x"00",	-- Hex Addr	7307	29447
x"00",	-- Hex Addr	7308	29448
x"00",	-- Hex Addr	7309	29449
x"00",	-- Hex Addr	730A	29450
x"00",	-- Hex Addr	730B	29451
x"00",	-- Hex Addr	730C	29452
x"00",	-- Hex Addr	730D	29453
x"00",	-- Hex Addr	730E	29454
x"00",	-- Hex Addr	730F	29455
x"00",	-- Hex Addr	7310	29456
x"00",	-- Hex Addr	7311	29457
x"00",	-- Hex Addr	7312	29458
x"00",	-- Hex Addr	7313	29459
x"00",	-- Hex Addr	7314	29460
x"00",	-- Hex Addr	7315	29461
x"00",	-- Hex Addr	7316	29462
x"00",	-- Hex Addr	7317	29463
x"00",	-- Hex Addr	7318	29464
x"00",	-- Hex Addr	7319	29465
x"00",	-- Hex Addr	731A	29466
x"00",	-- Hex Addr	731B	29467
x"00",	-- Hex Addr	731C	29468
x"00",	-- Hex Addr	731D	29469
x"00",	-- Hex Addr	731E	29470
x"00",	-- Hex Addr	731F	29471
x"00",	-- Hex Addr	7320	29472
x"00",	-- Hex Addr	7321	29473
x"00",	-- Hex Addr	7322	29474
x"00",	-- Hex Addr	7323	29475
x"00",	-- Hex Addr	7324	29476
x"00",	-- Hex Addr	7325	29477
x"00",	-- Hex Addr	7326	29478
x"00",	-- Hex Addr	7327	29479
x"00",	-- Hex Addr	7328	29480
x"00",	-- Hex Addr	7329	29481
x"00",	-- Hex Addr	732A	29482
x"00",	-- Hex Addr	732B	29483
x"00",	-- Hex Addr	732C	29484
x"00",	-- Hex Addr	732D	29485
x"00",	-- Hex Addr	732E	29486
x"00",	-- Hex Addr	732F	29487
x"00",	-- Hex Addr	7330	29488
x"00",	-- Hex Addr	7331	29489
x"00",	-- Hex Addr	7332	29490
x"00",	-- Hex Addr	7333	29491
x"00",	-- Hex Addr	7334	29492
x"00",	-- Hex Addr	7335	29493
x"00",	-- Hex Addr	7336	29494
x"00",	-- Hex Addr	7337	29495
x"00",	-- Hex Addr	7338	29496
x"00",	-- Hex Addr	7339	29497
x"00",	-- Hex Addr	733A	29498
x"00",	-- Hex Addr	733B	29499
x"00",	-- Hex Addr	733C	29500
x"00",	-- Hex Addr	733D	29501
x"00",	-- Hex Addr	733E	29502
x"00",	-- Hex Addr	733F	29503
x"00",	-- Hex Addr	7340	29504
x"00",	-- Hex Addr	7341	29505
x"00",	-- Hex Addr	7342	29506
x"00",	-- Hex Addr	7343	29507
x"00",	-- Hex Addr	7344	29508
x"00",	-- Hex Addr	7345	29509
x"00",	-- Hex Addr	7346	29510
x"00",	-- Hex Addr	7347	29511
x"00",	-- Hex Addr	7348	29512
x"00",	-- Hex Addr	7349	29513
x"00",	-- Hex Addr	734A	29514
x"00",	-- Hex Addr	734B	29515
x"00",	-- Hex Addr	734C	29516
x"00",	-- Hex Addr	734D	29517
x"00",	-- Hex Addr	734E	29518
x"00",	-- Hex Addr	734F	29519
x"00",	-- Hex Addr	7350	29520
x"00",	-- Hex Addr	7351	29521
x"00",	-- Hex Addr	7352	29522
x"00",	-- Hex Addr	7353	29523
x"00",	-- Hex Addr	7354	29524
x"00",	-- Hex Addr	7355	29525
x"00",	-- Hex Addr	7356	29526
x"00",	-- Hex Addr	7357	29527
x"00",	-- Hex Addr	7358	29528
x"00",	-- Hex Addr	7359	29529
x"00",	-- Hex Addr	735A	29530
x"00",	-- Hex Addr	735B	29531
x"00",	-- Hex Addr	735C	29532
x"00",	-- Hex Addr	735D	29533
x"00",	-- Hex Addr	735E	29534
x"00",	-- Hex Addr	735F	29535
x"00",	-- Hex Addr	7360	29536
x"00",	-- Hex Addr	7361	29537
x"00",	-- Hex Addr	7362	29538
x"00",	-- Hex Addr	7363	29539
x"00",	-- Hex Addr	7364	29540
x"00",	-- Hex Addr	7365	29541
x"00",	-- Hex Addr	7366	29542
x"00",	-- Hex Addr	7367	29543
x"00",	-- Hex Addr	7368	29544
x"00",	-- Hex Addr	7369	29545
x"00",	-- Hex Addr	736A	29546
x"00",	-- Hex Addr	736B	29547
x"00",	-- Hex Addr	736C	29548
x"00",	-- Hex Addr	736D	29549
x"00",	-- Hex Addr	736E	29550
x"00",	-- Hex Addr	736F	29551
x"00",	-- Hex Addr	7370	29552
x"00",	-- Hex Addr	7371	29553
x"00",	-- Hex Addr	7372	29554
x"00",	-- Hex Addr	7373	29555
x"00",	-- Hex Addr	7374	29556
x"00",	-- Hex Addr	7375	29557
x"00",	-- Hex Addr	7376	29558
x"00",	-- Hex Addr	7377	29559
x"00",	-- Hex Addr	7378	29560
x"00",	-- Hex Addr	7379	29561
x"00",	-- Hex Addr	737A	29562
x"00",	-- Hex Addr	737B	29563
x"00",	-- Hex Addr	737C	29564
x"00",	-- Hex Addr	737D	29565
x"00",	-- Hex Addr	737E	29566
x"00",	-- Hex Addr	737F	29567
x"00",	-- Hex Addr	7380	29568
x"00",	-- Hex Addr	7381	29569
x"00",	-- Hex Addr	7382	29570
x"00",	-- Hex Addr	7383	29571
x"00",	-- Hex Addr	7384	29572
x"00",	-- Hex Addr	7385	29573
x"00",	-- Hex Addr	7386	29574
x"00",	-- Hex Addr	7387	29575
x"00",	-- Hex Addr	7388	29576
x"00",	-- Hex Addr	7389	29577
x"00",	-- Hex Addr	738A	29578
x"00",	-- Hex Addr	738B	29579
x"00",	-- Hex Addr	738C	29580
x"00",	-- Hex Addr	738D	29581
x"00",	-- Hex Addr	738E	29582
x"00",	-- Hex Addr	738F	29583
x"00",	-- Hex Addr	7390	29584
x"00",	-- Hex Addr	7391	29585
x"00",	-- Hex Addr	7392	29586
x"00",	-- Hex Addr	7393	29587
x"00",	-- Hex Addr	7394	29588
x"00",	-- Hex Addr	7395	29589
x"00",	-- Hex Addr	7396	29590
x"00",	-- Hex Addr	7397	29591
x"00",	-- Hex Addr	7398	29592
x"00",	-- Hex Addr	7399	29593
x"00",	-- Hex Addr	739A	29594
x"00",	-- Hex Addr	739B	29595
x"00",	-- Hex Addr	739C	29596
x"00",	-- Hex Addr	739D	29597
x"00",	-- Hex Addr	739E	29598
x"00",	-- Hex Addr	739F	29599
x"00",	-- Hex Addr	73A0	29600
x"00",	-- Hex Addr	73A1	29601
x"00",	-- Hex Addr	73A2	29602
x"00",	-- Hex Addr	73A3	29603
x"00",	-- Hex Addr	73A4	29604
x"00",	-- Hex Addr	73A5	29605
x"00",	-- Hex Addr	73A6	29606
x"00",	-- Hex Addr	73A7	29607
x"00",	-- Hex Addr	73A8	29608
x"00",	-- Hex Addr	73A9	29609
x"00",	-- Hex Addr	73AA	29610
x"00",	-- Hex Addr	73AB	29611
x"00",	-- Hex Addr	73AC	29612
x"00",	-- Hex Addr	73AD	29613
x"00",	-- Hex Addr	73AE	29614
x"00",	-- Hex Addr	73AF	29615
x"00",	-- Hex Addr	73B0	29616
x"00",	-- Hex Addr	73B1	29617
x"00",	-- Hex Addr	73B2	29618
x"00",	-- Hex Addr	73B3	29619
x"00",	-- Hex Addr	73B4	29620
x"00",	-- Hex Addr	73B5	29621
x"00",	-- Hex Addr	73B6	29622
x"00",	-- Hex Addr	73B7	29623
x"00",	-- Hex Addr	73B8	29624
x"00",	-- Hex Addr	73B9	29625
x"00",	-- Hex Addr	73BA	29626
x"00",	-- Hex Addr	73BB	29627
x"00",	-- Hex Addr	73BC	29628
x"00",	-- Hex Addr	73BD	29629
x"00",	-- Hex Addr	73BE	29630
x"00",	-- Hex Addr	73BF	29631
x"00",	-- Hex Addr	73C0	29632
x"00",	-- Hex Addr	73C1	29633
x"00",	-- Hex Addr	73C2	29634
x"00",	-- Hex Addr	73C3	29635
x"00",	-- Hex Addr	73C4	29636
x"00",	-- Hex Addr	73C5	29637
x"00",	-- Hex Addr	73C6	29638
x"00",	-- Hex Addr	73C7	29639
x"00",	-- Hex Addr	73C8	29640
x"00",	-- Hex Addr	73C9	29641
x"00",	-- Hex Addr	73CA	29642
x"00",	-- Hex Addr	73CB	29643
x"00",	-- Hex Addr	73CC	29644
x"00",	-- Hex Addr	73CD	29645
x"00",	-- Hex Addr	73CE	29646
x"00",	-- Hex Addr	73CF	29647
x"00",	-- Hex Addr	73D0	29648
x"00",	-- Hex Addr	73D1	29649
x"00",	-- Hex Addr	73D2	29650
x"00",	-- Hex Addr	73D3	29651
x"00",	-- Hex Addr	73D4	29652
x"00",	-- Hex Addr	73D5	29653
x"00",	-- Hex Addr	73D6	29654
x"00",	-- Hex Addr	73D7	29655
x"00",	-- Hex Addr	73D8	29656
x"00",	-- Hex Addr	73D9	29657
x"00",	-- Hex Addr	73DA	29658
x"00",	-- Hex Addr	73DB	29659
x"00",	-- Hex Addr	73DC	29660
x"00",	-- Hex Addr	73DD	29661
x"00",	-- Hex Addr	73DE	29662
x"00",	-- Hex Addr	73DF	29663
x"00",	-- Hex Addr	73E0	29664
x"00",	-- Hex Addr	73E1	29665
x"00",	-- Hex Addr	73E2	29666
x"00",	-- Hex Addr	73E3	29667
x"00",	-- Hex Addr	73E4	29668
x"00",	-- Hex Addr	73E5	29669
x"00",	-- Hex Addr	73E6	29670
x"00",	-- Hex Addr	73E7	29671
x"00",	-- Hex Addr	73E8	29672
x"00",	-- Hex Addr	73E9	29673
x"00",	-- Hex Addr	73EA	29674
x"00",	-- Hex Addr	73EB	29675
x"00",	-- Hex Addr	73EC	29676
x"00",	-- Hex Addr	73ED	29677
x"00",	-- Hex Addr	73EE	29678
x"00",	-- Hex Addr	73EF	29679
x"00",	-- Hex Addr	73F0	29680
x"00",	-- Hex Addr	73F1	29681
x"00",	-- Hex Addr	73F2	29682
x"00",	-- Hex Addr	73F3	29683
x"00",	-- Hex Addr	73F4	29684
x"00",	-- Hex Addr	73F5	29685
x"00",	-- Hex Addr	73F6	29686
x"00",	-- Hex Addr	73F7	29687
x"00",	-- Hex Addr	73F8	29688
x"00",	-- Hex Addr	73F9	29689
x"00",	-- Hex Addr	73FA	29690
x"00",	-- Hex Addr	73FB	29691
x"00",	-- Hex Addr	73FC	29692
x"00",	-- Hex Addr	73FD	29693
x"00",	-- Hex Addr	73FE	29694
x"00",	-- Hex Addr	73FF	29695
x"00",	-- Hex Addr	7400	29696
x"00",	-- Hex Addr	7401	29697
x"00",	-- Hex Addr	7402	29698
x"00",	-- Hex Addr	7403	29699
x"00",	-- Hex Addr	7404	29700
x"00",	-- Hex Addr	7405	29701
x"00",	-- Hex Addr	7406	29702
x"00",	-- Hex Addr	7407	29703
x"00",	-- Hex Addr	7408	29704
x"00",	-- Hex Addr	7409	29705
x"00",	-- Hex Addr	740A	29706
x"00",	-- Hex Addr	740B	29707
x"00",	-- Hex Addr	740C	29708
x"00",	-- Hex Addr	740D	29709
x"00",	-- Hex Addr	740E	29710
x"00",	-- Hex Addr	740F	29711
x"00",	-- Hex Addr	7410	29712
x"00",	-- Hex Addr	7411	29713
x"00",	-- Hex Addr	7412	29714
x"00",	-- Hex Addr	7413	29715
x"00",	-- Hex Addr	7414	29716
x"00",	-- Hex Addr	7415	29717
x"00",	-- Hex Addr	7416	29718
x"00",	-- Hex Addr	7417	29719
x"00",	-- Hex Addr	7418	29720
x"00",	-- Hex Addr	7419	29721
x"00",	-- Hex Addr	741A	29722
x"00",	-- Hex Addr	741B	29723
x"00",	-- Hex Addr	741C	29724
x"00",	-- Hex Addr	741D	29725
x"00",	-- Hex Addr	741E	29726
x"00",	-- Hex Addr	741F	29727
x"00",	-- Hex Addr	7420	29728
x"00",	-- Hex Addr	7421	29729
x"00",	-- Hex Addr	7422	29730
x"00",	-- Hex Addr	7423	29731
x"00",	-- Hex Addr	7424	29732
x"00",	-- Hex Addr	7425	29733
x"00",	-- Hex Addr	7426	29734
x"00",	-- Hex Addr	7427	29735
x"00",	-- Hex Addr	7428	29736
x"00",	-- Hex Addr	7429	29737
x"00",	-- Hex Addr	742A	29738
x"00",	-- Hex Addr	742B	29739
x"00",	-- Hex Addr	742C	29740
x"00",	-- Hex Addr	742D	29741
x"00",	-- Hex Addr	742E	29742
x"00",	-- Hex Addr	742F	29743
x"00",	-- Hex Addr	7430	29744
x"00",	-- Hex Addr	7431	29745
x"00",	-- Hex Addr	7432	29746
x"00",	-- Hex Addr	7433	29747
x"00",	-- Hex Addr	7434	29748
x"00",	-- Hex Addr	7435	29749
x"00",	-- Hex Addr	7436	29750
x"00",	-- Hex Addr	7437	29751
x"00",	-- Hex Addr	7438	29752
x"00",	-- Hex Addr	7439	29753
x"00",	-- Hex Addr	743A	29754
x"00",	-- Hex Addr	743B	29755
x"00",	-- Hex Addr	743C	29756
x"00",	-- Hex Addr	743D	29757
x"00",	-- Hex Addr	743E	29758
x"00",	-- Hex Addr	743F	29759
x"00",	-- Hex Addr	7440	29760
x"00",	-- Hex Addr	7441	29761
x"00",	-- Hex Addr	7442	29762
x"00",	-- Hex Addr	7443	29763
x"00",	-- Hex Addr	7444	29764
x"00",	-- Hex Addr	7445	29765
x"00",	-- Hex Addr	7446	29766
x"00",	-- Hex Addr	7447	29767
x"00",	-- Hex Addr	7448	29768
x"00",	-- Hex Addr	7449	29769
x"00",	-- Hex Addr	744A	29770
x"00",	-- Hex Addr	744B	29771
x"00",	-- Hex Addr	744C	29772
x"00",	-- Hex Addr	744D	29773
x"00",	-- Hex Addr	744E	29774
x"00",	-- Hex Addr	744F	29775
x"00",	-- Hex Addr	7450	29776
x"00",	-- Hex Addr	7451	29777
x"00",	-- Hex Addr	7452	29778
x"00",	-- Hex Addr	7453	29779
x"00",	-- Hex Addr	7454	29780
x"00",	-- Hex Addr	7455	29781
x"00",	-- Hex Addr	7456	29782
x"00",	-- Hex Addr	7457	29783
x"00",	-- Hex Addr	7458	29784
x"00",	-- Hex Addr	7459	29785
x"00",	-- Hex Addr	745A	29786
x"00",	-- Hex Addr	745B	29787
x"00",	-- Hex Addr	745C	29788
x"00",	-- Hex Addr	745D	29789
x"00",	-- Hex Addr	745E	29790
x"00",	-- Hex Addr	745F	29791
x"00",	-- Hex Addr	7460	29792
x"00",	-- Hex Addr	7461	29793
x"00",	-- Hex Addr	7462	29794
x"00",	-- Hex Addr	7463	29795
x"00",	-- Hex Addr	7464	29796
x"00",	-- Hex Addr	7465	29797
x"00",	-- Hex Addr	7466	29798
x"00",	-- Hex Addr	7467	29799
x"00",	-- Hex Addr	7468	29800
x"00",	-- Hex Addr	7469	29801
x"00",	-- Hex Addr	746A	29802
x"00",	-- Hex Addr	746B	29803
x"00",	-- Hex Addr	746C	29804
x"00",	-- Hex Addr	746D	29805
x"00",	-- Hex Addr	746E	29806
x"00",	-- Hex Addr	746F	29807
x"00",	-- Hex Addr	7470	29808
x"00",	-- Hex Addr	7471	29809
x"00",	-- Hex Addr	7472	29810
x"00",	-- Hex Addr	7473	29811
x"00",	-- Hex Addr	7474	29812
x"00",	-- Hex Addr	7475	29813
x"00",	-- Hex Addr	7476	29814
x"00",	-- Hex Addr	7477	29815
x"00",	-- Hex Addr	7478	29816
x"00",	-- Hex Addr	7479	29817
x"00",	-- Hex Addr	747A	29818
x"00",	-- Hex Addr	747B	29819
x"00",	-- Hex Addr	747C	29820
x"00",	-- Hex Addr	747D	29821
x"00",	-- Hex Addr	747E	29822
x"00",	-- Hex Addr	747F	29823
x"00",	-- Hex Addr	7480	29824
x"00",	-- Hex Addr	7481	29825
x"00",	-- Hex Addr	7482	29826
x"00",	-- Hex Addr	7483	29827
x"00",	-- Hex Addr	7484	29828
x"00",	-- Hex Addr	7485	29829
x"00",	-- Hex Addr	7486	29830
x"00",	-- Hex Addr	7487	29831
x"00",	-- Hex Addr	7488	29832
x"00",	-- Hex Addr	7489	29833
x"00",	-- Hex Addr	748A	29834
x"00",	-- Hex Addr	748B	29835
x"00",	-- Hex Addr	748C	29836
x"00",	-- Hex Addr	748D	29837
x"00",	-- Hex Addr	748E	29838
x"00",	-- Hex Addr	748F	29839
x"00",	-- Hex Addr	7490	29840
x"00",	-- Hex Addr	7491	29841
x"00",	-- Hex Addr	7492	29842
x"00",	-- Hex Addr	7493	29843
x"00",	-- Hex Addr	7494	29844
x"00",	-- Hex Addr	7495	29845
x"00",	-- Hex Addr	7496	29846
x"00",	-- Hex Addr	7497	29847
x"00",	-- Hex Addr	7498	29848
x"00",	-- Hex Addr	7499	29849
x"00",	-- Hex Addr	749A	29850
x"00",	-- Hex Addr	749B	29851
x"00",	-- Hex Addr	749C	29852
x"00",	-- Hex Addr	749D	29853
x"00",	-- Hex Addr	749E	29854
x"00",	-- Hex Addr	749F	29855
x"00",	-- Hex Addr	74A0	29856
x"00",	-- Hex Addr	74A1	29857
x"00",	-- Hex Addr	74A2	29858
x"00",	-- Hex Addr	74A3	29859
x"00",	-- Hex Addr	74A4	29860
x"00",	-- Hex Addr	74A5	29861
x"00",	-- Hex Addr	74A6	29862
x"00",	-- Hex Addr	74A7	29863
x"00",	-- Hex Addr	74A8	29864
x"00",	-- Hex Addr	74A9	29865
x"00",	-- Hex Addr	74AA	29866
x"00",	-- Hex Addr	74AB	29867
x"00",	-- Hex Addr	74AC	29868
x"00",	-- Hex Addr	74AD	29869
x"00",	-- Hex Addr	74AE	29870
x"00",	-- Hex Addr	74AF	29871
x"00",	-- Hex Addr	74B0	29872
x"00",	-- Hex Addr	74B1	29873
x"00",	-- Hex Addr	74B2	29874
x"00",	-- Hex Addr	74B3	29875
x"00",	-- Hex Addr	74B4	29876
x"00",	-- Hex Addr	74B5	29877
x"00",	-- Hex Addr	74B6	29878
x"00",	-- Hex Addr	74B7	29879
x"00",	-- Hex Addr	74B8	29880
x"00",	-- Hex Addr	74B9	29881
x"00",	-- Hex Addr	74BA	29882
x"00",	-- Hex Addr	74BB	29883
x"00",	-- Hex Addr	74BC	29884
x"00",	-- Hex Addr	74BD	29885
x"00",	-- Hex Addr	74BE	29886
x"00",	-- Hex Addr	74BF	29887
x"00",	-- Hex Addr	74C0	29888
x"00",	-- Hex Addr	74C1	29889
x"00",	-- Hex Addr	74C2	29890
x"00",	-- Hex Addr	74C3	29891
x"00",	-- Hex Addr	74C4	29892
x"00",	-- Hex Addr	74C5	29893
x"00",	-- Hex Addr	74C6	29894
x"00",	-- Hex Addr	74C7	29895
x"00",	-- Hex Addr	74C8	29896
x"00",	-- Hex Addr	74C9	29897
x"00",	-- Hex Addr	74CA	29898
x"00",	-- Hex Addr	74CB	29899
x"00",	-- Hex Addr	74CC	29900
x"00",	-- Hex Addr	74CD	29901
x"00",	-- Hex Addr	74CE	29902
x"00",	-- Hex Addr	74CF	29903
x"00",	-- Hex Addr	74D0	29904
x"00",	-- Hex Addr	74D1	29905
x"00",	-- Hex Addr	74D2	29906
x"00",	-- Hex Addr	74D3	29907
x"00",	-- Hex Addr	74D4	29908
x"00",	-- Hex Addr	74D5	29909
x"00",	-- Hex Addr	74D6	29910
x"00",	-- Hex Addr	74D7	29911
x"00",	-- Hex Addr	74D8	29912
x"00",	-- Hex Addr	74D9	29913
x"00",	-- Hex Addr	74DA	29914
x"00",	-- Hex Addr	74DB	29915
x"00",	-- Hex Addr	74DC	29916
x"00",	-- Hex Addr	74DD	29917
x"00",	-- Hex Addr	74DE	29918
x"00",	-- Hex Addr	74DF	29919
x"00",	-- Hex Addr	74E0	29920
x"00",	-- Hex Addr	74E1	29921
x"00",	-- Hex Addr	74E2	29922
x"00",	-- Hex Addr	74E3	29923
x"00",	-- Hex Addr	74E4	29924
x"00",	-- Hex Addr	74E5	29925
x"00",	-- Hex Addr	74E6	29926
x"00",	-- Hex Addr	74E7	29927
x"00",	-- Hex Addr	74E8	29928
x"00",	-- Hex Addr	74E9	29929
x"00",	-- Hex Addr	74EA	29930
x"00",	-- Hex Addr	74EB	29931
x"00",	-- Hex Addr	74EC	29932
x"00",	-- Hex Addr	74ED	29933
x"00",	-- Hex Addr	74EE	29934
x"00",	-- Hex Addr	74EF	29935
x"00",	-- Hex Addr	74F0	29936
x"00",	-- Hex Addr	74F1	29937
x"00",	-- Hex Addr	74F2	29938
x"00",	-- Hex Addr	74F3	29939
x"00",	-- Hex Addr	74F4	29940
x"00",	-- Hex Addr	74F5	29941
x"00",	-- Hex Addr	74F6	29942
x"00",	-- Hex Addr	74F7	29943
x"00",	-- Hex Addr	74F8	29944
x"00",	-- Hex Addr	74F9	29945
x"00",	-- Hex Addr	74FA	29946
x"00",	-- Hex Addr	74FB	29947
x"00",	-- Hex Addr	74FC	29948
x"00",	-- Hex Addr	74FD	29949
x"00",	-- Hex Addr	74FE	29950
x"00",	-- Hex Addr	74FF	29951
x"00",	-- Hex Addr	7500	29952
x"00",	-- Hex Addr	7501	29953
x"00",	-- Hex Addr	7502	29954
x"00",	-- Hex Addr	7503	29955
x"00",	-- Hex Addr	7504	29956
x"00",	-- Hex Addr	7505	29957
x"00",	-- Hex Addr	7506	29958
x"00",	-- Hex Addr	7507	29959
x"00",	-- Hex Addr	7508	29960
x"00",	-- Hex Addr	7509	29961
x"00",	-- Hex Addr	750A	29962
x"00",	-- Hex Addr	750B	29963
x"00",	-- Hex Addr	750C	29964
x"00",	-- Hex Addr	750D	29965
x"00",	-- Hex Addr	750E	29966
x"00",	-- Hex Addr	750F	29967
x"00",	-- Hex Addr	7510	29968
x"00",	-- Hex Addr	7511	29969
x"00",	-- Hex Addr	7512	29970
x"00",	-- Hex Addr	7513	29971
x"00",	-- Hex Addr	7514	29972
x"00",	-- Hex Addr	7515	29973
x"00",	-- Hex Addr	7516	29974
x"00",	-- Hex Addr	7517	29975
x"00",	-- Hex Addr	7518	29976
x"00",	-- Hex Addr	7519	29977
x"00",	-- Hex Addr	751A	29978
x"00",	-- Hex Addr	751B	29979
x"00",	-- Hex Addr	751C	29980
x"00",	-- Hex Addr	751D	29981
x"00",	-- Hex Addr	751E	29982
x"00",	-- Hex Addr	751F	29983
x"00",	-- Hex Addr	7520	29984
x"00",	-- Hex Addr	7521	29985
x"00",	-- Hex Addr	7522	29986
x"00",	-- Hex Addr	7523	29987
x"00",	-- Hex Addr	7524	29988
x"00",	-- Hex Addr	7525	29989
x"00",	-- Hex Addr	7526	29990
x"00",	-- Hex Addr	7527	29991
x"00",	-- Hex Addr	7528	29992
x"00",	-- Hex Addr	7529	29993
x"00",	-- Hex Addr	752A	29994
x"00",	-- Hex Addr	752B	29995
x"00",	-- Hex Addr	752C	29996
x"00",	-- Hex Addr	752D	29997
x"00",	-- Hex Addr	752E	29998
x"00",	-- Hex Addr	752F	29999
x"00",	-- Hex Addr	7530	30000
x"00",	-- Hex Addr	7531	30001
x"00",	-- Hex Addr	7532	30002
x"00",	-- Hex Addr	7533	30003
x"00",	-- Hex Addr	7534	30004
x"00",	-- Hex Addr	7535	30005
x"00",	-- Hex Addr	7536	30006
x"00",	-- Hex Addr	7537	30007
x"00",	-- Hex Addr	7538	30008
x"00",	-- Hex Addr	7539	30009
x"00",	-- Hex Addr	753A	30010
x"00",	-- Hex Addr	753B	30011
x"00",	-- Hex Addr	753C	30012
x"00",	-- Hex Addr	753D	30013
x"00",	-- Hex Addr	753E	30014
x"00",	-- Hex Addr	753F	30015
x"00",	-- Hex Addr	7540	30016
x"00",	-- Hex Addr	7541	30017
x"00",	-- Hex Addr	7542	30018
x"00",	-- Hex Addr	7543	30019
x"00",	-- Hex Addr	7544	30020
x"00",	-- Hex Addr	7545	30021
x"00",	-- Hex Addr	7546	30022
x"00",	-- Hex Addr	7547	30023
x"00",	-- Hex Addr	7548	30024
x"00",	-- Hex Addr	7549	30025
x"00",	-- Hex Addr	754A	30026
x"00",	-- Hex Addr	754B	30027
x"00",	-- Hex Addr	754C	30028
x"00",	-- Hex Addr	754D	30029
x"00",	-- Hex Addr	754E	30030
x"00",	-- Hex Addr	754F	30031
x"00",	-- Hex Addr	7550	30032
x"00",	-- Hex Addr	7551	30033
x"00",	-- Hex Addr	7552	30034
x"00",	-- Hex Addr	7553	30035
x"00",	-- Hex Addr	7554	30036
x"00",	-- Hex Addr	7555	30037
x"00",	-- Hex Addr	7556	30038
x"00",	-- Hex Addr	7557	30039
x"00",	-- Hex Addr	7558	30040
x"00",	-- Hex Addr	7559	30041
x"00",	-- Hex Addr	755A	30042
x"00",	-- Hex Addr	755B	30043
x"00",	-- Hex Addr	755C	30044
x"00",	-- Hex Addr	755D	30045
x"00",	-- Hex Addr	755E	30046
x"00",	-- Hex Addr	755F	30047
x"00",	-- Hex Addr	7560	30048
x"00",	-- Hex Addr	7561	30049
x"00",	-- Hex Addr	7562	30050
x"00",	-- Hex Addr	7563	30051
x"00",	-- Hex Addr	7564	30052
x"00",	-- Hex Addr	7565	30053
x"00",	-- Hex Addr	7566	30054
x"00",	-- Hex Addr	7567	30055
x"00",	-- Hex Addr	7568	30056
x"00",	-- Hex Addr	7569	30057
x"00",	-- Hex Addr	756A	30058
x"00",	-- Hex Addr	756B	30059
x"00",	-- Hex Addr	756C	30060
x"00",	-- Hex Addr	756D	30061
x"00",	-- Hex Addr	756E	30062
x"00",	-- Hex Addr	756F	30063
x"00",	-- Hex Addr	7570	30064
x"00",	-- Hex Addr	7571	30065
x"00",	-- Hex Addr	7572	30066
x"00",	-- Hex Addr	7573	30067
x"00",	-- Hex Addr	7574	30068
x"00",	-- Hex Addr	7575	30069
x"00",	-- Hex Addr	7576	30070
x"00",	-- Hex Addr	7577	30071
x"00",	-- Hex Addr	7578	30072
x"00",	-- Hex Addr	7579	30073
x"00",	-- Hex Addr	757A	30074
x"00",	-- Hex Addr	757B	30075
x"00",	-- Hex Addr	757C	30076
x"00",	-- Hex Addr	757D	30077
x"00",	-- Hex Addr	757E	30078
x"00",	-- Hex Addr	757F	30079
x"00",	-- Hex Addr	7580	30080
x"00",	-- Hex Addr	7581	30081
x"00",	-- Hex Addr	7582	30082
x"00",	-- Hex Addr	7583	30083
x"00",	-- Hex Addr	7584	30084
x"00",	-- Hex Addr	7585	30085
x"00",	-- Hex Addr	7586	30086
x"00",	-- Hex Addr	7587	30087
x"00",	-- Hex Addr	7588	30088
x"00",	-- Hex Addr	7589	30089
x"00",	-- Hex Addr	758A	30090
x"00",	-- Hex Addr	758B	30091
x"00",	-- Hex Addr	758C	30092
x"00",	-- Hex Addr	758D	30093
x"00",	-- Hex Addr	758E	30094
x"00",	-- Hex Addr	758F	30095
x"00",	-- Hex Addr	7590	30096
x"00",	-- Hex Addr	7591	30097
x"00",	-- Hex Addr	7592	30098
x"00",	-- Hex Addr	7593	30099
x"00",	-- Hex Addr	7594	30100
x"00",	-- Hex Addr	7595	30101
x"00",	-- Hex Addr	7596	30102
x"00",	-- Hex Addr	7597	30103
x"00",	-- Hex Addr	7598	30104
x"00",	-- Hex Addr	7599	30105
x"00",	-- Hex Addr	759A	30106
x"00",	-- Hex Addr	759B	30107
x"00",	-- Hex Addr	759C	30108
x"00",	-- Hex Addr	759D	30109
x"00",	-- Hex Addr	759E	30110
x"00",	-- Hex Addr	759F	30111
x"00",	-- Hex Addr	75A0	30112
x"00",	-- Hex Addr	75A1	30113
x"00",	-- Hex Addr	75A2	30114
x"00",	-- Hex Addr	75A3	30115
x"00",	-- Hex Addr	75A4	30116
x"00",	-- Hex Addr	75A5	30117
x"00",	-- Hex Addr	75A6	30118
x"00",	-- Hex Addr	75A7	30119
x"00",	-- Hex Addr	75A8	30120
x"00",	-- Hex Addr	75A9	30121
x"00",	-- Hex Addr	75AA	30122
x"00",	-- Hex Addr	75AB	30123
x"00",	-- Hex Addr	75AC	30124
x"00",	-- Hex Addr	75AD	30125
x"00",	-- Hex Addr	75AE	30126
x"00",	-- Hex Addr	75AF	30127
x"00",	-- Hex Addr	75B0	30128
x"00",	-- Hex Addr	75B1	30129
x"00",	-- Hex Addr	75B2	30130
x"00",	-- Hex Addr	75B3	30131
x"00",	-- Hex Addr	75B4	30132
x"00",	-- Hex Addr	75B5	30133
x"00",	-- Hex Addr	75B6	30134
x"00",	-- Hex Addr	75B7	30135
x"00",	-- Hex Addr	75B8	30136
x"00",	-- Hex Addr	75B9	30137
x"00",	-- Hex Addr	75BA	30138
x"00",	-- Hex Addr	75BB	30139
x"00",	-- Hex Addr	75BC	30140
x"00",	-- Hex Addr	75BD	30141
x"00",	-- Hex Addr	75BE	30142
x"00",	-- Hex Addr	75BF	30143
x"00",	-- Hex Addr	75C0	30144
x"00",	-- Hex Addr	75C1	30145
x"00",	-- Hex Addr	75C2	30146
x"00",	-- Hex Addr	75C3	30147
x"00",	-- Hex Addr	75C4	30148
x"00",	-- Hex Addr	75C5	30149
x"00",	-- Hex Addr	75C6	30150
x"00",	-- Hex Addr	75C7	30151
x"00",	-- Hex Addr	75C8	30152
x"00",	-- Hex Addr	75C9	30153
x"00",	-- Hex Addr	75CA	30154
x"00",	-- Hex Addr	75CB	30155
x"00",	-- Hex Addr	75CC	30156
x"00",	-- Hex Addr	75CD	30157
x"00",	-- Hex Addr	75CE	30158
x"00",	-- Hex Addr	75CF	30159
x"00",	-- Hex Addr	75D0	30160
x"00",	-- Hex Addr	75D1	30161
x"00",	-- Hex Addr	75D2	30162
x"00",	-- Hex Addr	75D3	30163
x"00",	-- Hex Addr	75D4	30164
x"00",	-- Hex Addr	75D5	30165
x"00",	-- Hex Addr	75D6	30166
x"00",	-- Hex Addr	75D7	30167
x"00",	-- Hex Addr	75D8	30168
x"00",	-- Hex Addr	75D9	30169
x"00",	-- Hex Addr	75DA	30170
x"00",	-- Hex Addr	75DB	30171
x"00",	-- Hex Addr	75DC	30172
x"00",	-- Hex Addr	75DD	30173
x"00",	-- Hex Addr	75DE	30174
x"00",	-- Hex Addr	75DF	30175
x"00",	-- Hex Addr	75E0	30176
x"00",	-- Hex Addr	75E1	30177
x"00",	-- Hex Addr	75E2	30178
x"00",	-- Hex Addr	75E3	30179
x"00",	-- Hex Addr	75E4	30180
x"00",	-- Hex Addr	75E5	30181
x"00",	-- Hex Addr	75E6	30182
x"00",	-- Hex Addr	75E7	30183
x"00",	-- Hex Addr	75E8	30184
x"00",	-- Hex Addr	75E9	30185
x"00",	-- Hex Addr	75EA	30186
x"00",	-- Hex Addr	75EB	30187
x"00",	-- Hex Addr	75EC	30188
x"00",	-- Hex Addr	75ED	30189
x"00",	-- Hex Addr	75EE	30190
x"00",	-- Hex Addr	75EF	30191
x"00",	-- Hex Addr	75F0	30192
x"00",	-- Hex Addr	75F1	30193
x"00",	-- Hex Addr	75F2	30194
x"00",	-- Hex Addr	75F3	30195
x"00",	-- Hex Addr	75F4	30196
x"00",	-- Hex Addr	75F5	30197
x"00",	-- Hex Addr	75F6	30198
x"00",	-- Hex Addr	75F7	30199
x"00",	-- Hex Addr	75F8	30200
x"00",	-- Hex Addr	75F9	30201
x"00",	-- Hex Addr	75FA	30202
x"00",	-- Hex Addr	75FB	30203
x"00",	-- Hex Addr	75FC	30204
x"00",	-- Hex Addr	75FD	30205
x"00",	-- Hex Addr	75FE	30206
x"00",	-- Hex Addr	75FF	30207
x"00",	-- Hex Addr	7600	30208
x"00",	-- Hex Addr	7601	30209
x"00",	-- Hex Addr	7602	30210
x"00",	-- Hex Addr	7603	30211
x"00",	-- Hex Addr	7604	30212
x"00",	-- Hex Addr	7605	30213
x"00",	-- Hex Addr	7606	30214
x"00",	-- Hex Addr	7607	30215
x"00",	-- Hex Addr	7608	30216
x"00",	-- Hex Addr	7609	30217
x"00",	-- Hex Addr	760A	30218
x"00",	-- Hex Addr	760B	30219
x"00",	-- Hex Addr	760C	30220
x"00",	-- Hex Addr	760D	30221
x"00",	-- Hex Addr	760E	30222
x"00",	-- Hex Addr	760F	30223
x"00",	-- Hex Addr	7610	30224
x"00",	-- Hex Addr	7611	30225
x"00",	-- Hex Addr	7612	30226
x"00",	-- Hex Addr	7613	30227
x"00",	-- Hex Addr	7614	30228
x"00",	-- Hex Addr	7615	30229
x"00",	-- Hex Addr	7616	30230
x"00",	-- Hex Addr	7617	30231
x"00",	-- Hex Addr	7618	30232
x"00",	-- Hex Addr	7619	30233
x"00",	-- Hex Addr	761A	30234
x"00",	-- Hex Addr	761B	30235
x"00",	-- Hex Addr	761C	30236
x"00",	-- Hex Addr	761D	30237
x"00",	-- Hex Addr	761E	30238
x"00",	-- Hex Addr	761F	30239
x"00",	-- Hex Addr	7620	30240
x"00",	-- Hex Addr	7621	30241
x"00",	-- Hex Addr	7622	30242
x"00",	-- Hex Addr	7623	30243
x"00",	-- Hex Addr	7624	30244
x"00",	-- Hex Addr	7625	30245
x"00",	-- Hex Addr	7626	30246
x"00",	-- Hex Addr	7627	30247
x"00",	-- Hex Addr	7628	30248
x"00",	-- Hex Addr	7629	30249
x"00",	-- Hex Addr	762A	30250
x"00",	-- Hex Addr	762B	30251
x"00",	-- Hex Addr	762C	30252
x"00",	-- Hex Addr	762D	30253
x"00",	-- Hex Addr	762E	30254
x"00",	-- Hex Addr	762F	30255
x"00",	-- Hex Addr	7630	30256
x"00",	-- Hex Addr	7631	30257
x"00",	-- Hex Addr	7632	30258
x"00",	-- Hex Addr	7633	30259
x"00",	-- Hex Addr	7634	30260
x"00",	-- Hex Addr	7635	30261
x"00",	-- Hex Addr	7636	30262
x"00",	-- Hex Addr	7637	30263
x"00",	-- Hex Addr	7638	30264
x"00",	-- Hex Addr	7639	30265
x"00",	-- Hex Addr	763A	30266
x"00",	-- Hex Addr	763B	30267
x"00",	-- Hex Addr	763C	30268
x"00",	-- Hex Addr	763D	30269
x"00",	-- Hex Addr	763E	30270
x"00",	-- Hex Addr	763F	30271
x"00",	-- Hex Addr	7640	30272
x"00",	-- Hex Addr	7641	30273
x"00",	-- Hex Addr	7642	30274
x"00",	-- Hex Addr	7643	30275
x"00",	-- Hex Addr	7644	30276
x"00",	-- Hex Addr	7645	30277
x"00",	-- Hex Addr	7646	30278
x"00",	-- Hex Addr	7647	30279
x"00",	-- Hex Addr	7648	30280
x"00",	-- Hex Addr	7649	30281
x"00",	-- Hex Addr	764A	30282
x"00",	-- Hex Addr	764B	30283
x"00",	-- Hex Addr	764C	30284
x"00",	-- Hex Addr	764D	30285
x"00",	-- Hex Addr	764E	30286
x"00",	-- Hex Addr	764F	30287
x"00",	-- Hex Addr	7650	30288
x"00",	-- Hex Addr	7651	30289
x"00",	-- Hex Addr	7652	30290
x"00",	-- Hex Addr	7653	30291
x"00",	-- Hex Addr	7654	30292
x"00",	-- Hex Addr	7655	30293
x"00",	-- Hex Addr	7656	30294
x"00",	-- Hex Addr	7657	30295
x"00",	-- Hex Addr	7658	30296
x"00",	-- Hex Addr	7659	30297
x"00",	-- Hex Addr	765A	30298
x"00",	-- Hex Addr	765B	30299
x"00",	-- Hex Addr	765C	30300
x"00",	-- Hex Addr	765D	30301
x"00",	-- Hex Addr	765E	30302
x"00",	-- Hex Addr	765F	30303
x"00",	-- Hex Addr	7660	30304
x"00",	-- Hex Addr	7661	30305
x"00",	-- Hex Addr	7662	30306
x"00",	-- Hex Addr	7663	30307
x"00",	-- Hex Addr	7664	30308
x"00",	-- Hex Addr	7665	30309
x"00",	-- Hex Addr	7666	30310
x"00",	-- Hex Addr	7667	30311
x"00",	-- Hex Addr	7668	30312
x"00",	-- Hex Addr	7669	30313
x"00",	-- Hex Addr	766A	30314
x"00",	-- Hex Addr	766B	30315
x"00",	-- Hex Addr	766C	30316
x"00",	-- Hex Addr	766D	30317
x"00",	-- Hex Addr	766E	30318
x"00",	-- Hex Addr	766F	30319
x"00",	-- Hex Addr	7670	30320
x"00",	-- Hex Addr	7671	30321
x"00",	-- Hex Addr	7672	30322
x"00",	-- Hex Addr	7673	30323
x"00",	-- Hex Addr	7674	30324
x"00",	-- Hex Addr	7675	30325
x"00",	-- Hex Addr	7676	30326
x"00",	-- Hex Addr	7677	30327
x"00",	-- Hex Addr	7678	30328
x"00",	-- Hex Addr	7679	30329
x"00",	-- Hex Addr	767A	30330
x"00",	-- Hex Addr	767B	30331
x"00",	-- Hex Addr	767C	30332
x"00",	-- Hex Addr	767D	30333
x"00",	-- Hex Addr	767E	30334
x"00",	-- Hex Addr	767F	30335
x"00",	-- Hex Addr	7680	30336
x"00",	-- Hex Addr	7681	30337
x"00",	-- Hex Addr	7682	30338
x"00",	-- Hex Addr	7683	30339
x"00",	-- Hex Addr	7684	30340
x"00",	-- Hex Addr	7685	30341
x"00",	-- Hex Addr	7686	30342
x"00",	-- Hex Addr	7687	30343
x"00",	-- Hex Addr	7688	30344
x"00",	-- Hex Addr	7689	30345
x"00",	-- Hex Addr	768A	30346
x"00",	-- Hex Addr	768B	30347
x"00",	-- Hex Addr	768C	30348
x"00",	-- Hex Addr	768D	30349
x"00",	-- Hex Addr	768E	30350
x"00",	-- Hex Addr	768F	30351
x"00",	-- Hex Addr	7690	30352
x"00",	-- Hex Addr	7691	30353
x"00",	-- Hex Addr	7692	30354
x"00",	-- Hex Addr	7693	30355
x"00",	-- Hex Addr	7694	30356
x"00",	-- Hex Addr	7695	30357
x"00",	-- Hex Addr	7696	30358
x"00",	-- Hex Addr	7697	30359
x"00",	-- Hex Addr	7698	30360
x"00",	-- Hex Addr	7699	30361
x"00",	-- Hex Addr	769A	30362
x"00",	-- Hex Addr	769B	30363
x"00",	-- Hex Addr	769C	30364
x"00",	-- Hex Addr	769D	30365
x"00",	-- Hex Addr	769E	30366
x"00",	-- Hex Addr	769F	30367
x"00",	-- Hex Addr	76A0	30368
x"00",	-- Hex Addr	76A1	30369
x"00",	-- Hex Addr	76A2	30370
x"00",	-- Hex Addr	76A3	30371
x"00",	-- Hex Addr	76A4	30372
x"00",	-- Hex Addr	76A5	30373
x"00",	-- Hex Addr	76A6	30374
x"00",	-- Hex Addr	76A7	30375
x"00",	-- Hex Addr	76A8	30376
x"00",	-- Hex Addr	76A9	30377
x"00",	-- Hex Addr	76AA	30378
x"00",	-- Hex Addr	76AB	30379
x"00",	-- Hex Addr	76AC	30380
x"00",	-- Hex Addr	76AD	30381
x"00",	-- Hex Addr	76AE	30382
x"00",	-- Hex Addr	76AF	30383
x"00",	-- Hex Addr	76B0	30384
x"00",	-- Hex Addr	76B1	30385
x"00",	-- Hex Addr	76B2	30386
x"00",	-- Hex Addr	76B3	30387
x"00",	-- Hex Addr	76B4	30388
x"00",	-- Hex Addr	76B5	30389
x"00",	-- Hex Addr	76B6	30390
x"00",	-- Hex Addr	76B7	30391
x"00",	-- Hex Addr	76B8	30392
x"00",	-- Hex Addr	76B9	30393
x"00",	-- Hex Addr	76BA	30394
x"00",	-- Hex Addr	76BB	30395
x"00",	-- Hex Addr	76BC	30396
x"00",	-- Hex Addr	76BD	30397
x"00",	-- Hex Addr	76BE	30398
x"00",	-- Hex Addr	76BF	30399
x"00",	-- Hex Addr	76C0	30400
x"00",	-- Hex Addr	76C1	30401
x"00",	-- Hex Addr	76C2	30402
x"00",	-- Hex Addr	76C3	30403
x"00",	-- Hex Addr	76C4	30404
x"00",	-- Hex Addr	76C5	30405
x"00",	-- Hex Addr	76C6	30406
x"00",	-- Hex Addr	76C7	30407
x"00",	-- Hex Addr	76C8	30408
x"00",	-- Hex Addr	76C9	30409
x"00",	-- Hex Addr	76CA	30410
x"00",	-- Hex Addr	76CB	30411
x"00",	-- Hex Addr	76CC	30412
x"00",	-- Hex Addr	76CD	30413
x"00",	-- Hex Addr	76CE	30414
x"00",	-- Hex Addr	76CF	30415
x"00",	-- Hex Addr	76D0	30416
x"00",	-- Hex Addr	76D1	30417
x"00",	-- Hex Addr	76D2	30418
x"00",	-- Hex Addr	76D3	30419
x"00",	-- Hex Addr	76D4	30420
x"00",	-- Hex Addr	76D5	30421
x"00",	-- Hex Addr	76D6	30422
x"00",	-- Hex Addr	76D7	30423
x"00",	-- Hex Addr	76D8	30424
x"00",	-- Hex Addr	76D9	30425
x"00",	-- Hex Addr	76DA	30426
x"00",	-- Hex Addr	76DB	30427
x"00",	-- Hex Addr	76DC	30428
x"00",	-- Hex Addr	76DD	30429
x"00",	-- Hex Addr	76DE	30430
x"00",	-- Hex Addr	76DF	30431
x"00",	-- Hex Addr	76E0	30432
x"00",	-- Hex Addr	76E1	30433
x"00",	-- Hex Addr	76E2	30434
x"00",	-- Hex Addr	76E3	30435
x"00",	-- Hex Addr	76E4	30436
x"00",	-- Hex Addr	76E5	30437
x"00",	-- Hex Addr	76E6	30438
x"00",	-- Hex Addr	76E7	30439
x"00",	-- Hex Addr	76E8	30440
x"00",	-- Hex Addr	76E9	30441
x"00",	-- Hex Addr	76EA	30442
x"00",	-- Hex Addr	76EB	30443
x"00",	-- Hex Addr	76EC	30444
x"00",	-- Hex Addr	76ED	30445
x"00",	-- Hex Addr	76EE	30446
x"00",	-- Hex Addr	76EF	30447
x"00",	-- Hex Addr	76F0	30448
x"00",	-- Hex Addr	76F1	30449
x"00",	-- Hex Addr	76F2	30450
x"00",	-- Hex Addr	76F3	30451
x"00",	-- Hex Addr	76F4	30452
x"00",	-- Hex Addr	76F5	30453
x"00",	-- Hex Addr	76F6	30454
x"00",	-- Hex Addr	76F7	30455
x"00",	-- Hex Addr	76F8	30456
x"00",	-- Hex Addr	76F9	30457
x"00",	-- Hex Addr	76FA	30458
x"00",	-- Hex Addr	76FB	30459
x"00",	-- Hex Addr	76FC	30460
x"00",	-- Hex Addr	76FD	30461
x"00",	-- Hex Addr	76FE	30462
x"00",	-- Hex Addr	76FF	30463
x"00",	-- Hex Addr	7700	30464
x"00",	-- Hex Addr	7701	30465
x"00",	-- Hex Addr	7702	30466
x"00",	-- Hex Addr	7703	30467
x"00",	-- Hex Addr	7704	30468
x"00",	-- Hex Addr	7705	30469
x"00",	-- Hex Addr	7706	30470
x"00",	-- Hex Addr	7707	30471
x"00",	-- Hex Addr	7708	30472
x"00",	-- Hex Addr	7709	30473
x"00",	-- Hex Addr	770A	30474
x"00",	-- Hex Addr	770B	30475
x"00",	-- Hex Addr	770C	30476
x"00",	-- Hex Addr	770D	30477
x"00",	-- Hex Addr	770E	30478
x"00",	-- Hex Addr	770F	30479
x"00",	-- Hex Addr	7710	30480
x"00",	-- Hex Addr	7711	30481
x"00",	-- Hex Addr	7712	30482
x"00",	-- Hex Addr	7713	30483
x"00",	-- Hex Addr	7714	30484
x"00",	-- Hex Addr	7715	30485
x"00",	-- Hex Addr	7716	30486
x"00",	-- Hex Addr	7717	30487
x"00",	-- Hex Addr	7718	30488
x"00",	-- Hex Addr	7719	30489
x"00",	-- Hex Addr	771A	30490
x"00",	-- Hex Addr	771B	30491
x"00",	-- Hex Addr	771C	30492
x"00",	-- Hex Addr	771D	30493
x"00",	-- Hex Addr	771E	30494
x"00",	-- Hex Addr	771F	30495
x"00",	-- Hex Addr	7720	30496
x"00",	-- Hex Addr	7721	30497
x"00",	-- Hex Addr	7722	30498
x"00",	-- Hex Addr	7723	30499
x"00",	-- Hex Addr	7724	30500
x"00",	-- Hex Addr	7725	30501
x"00",	-- Hex Addr	7726	30502
x"00",	-- Hex Addr	7727	30503
x"00",	-- Hex Addr	7728	30504
x"00",	-- Hex Addr	7729	30505
x"00",	-- Hex Addr	772A	30506
x"00",	-- Hex Addr	772B	30507
x"00",	-- Hex Addr	772C	30508
x"00",	-- Hex Addr	772D	30509
x"00",	-- Hex Addr	772E	30510
x"00",	-- Hex Addr	772F	30511
x"00",	-- Hex Addr	7730	30512
x"00",	-- Hex Addr	7731	30513
x"00",	-- Hex Addr	7732	30514
x"00",	-- Hex Addr	7733	30515
x"00",	-- Hex Addr	7734	30516
x"00",	-- Hex Addr	7735	30517
x"00",	-- Hex Addr	7736	30518
x"00",	-- Hex Addr	7737	30519
x"00",	-- Hex Addr	7738	30520
x"00",	-- Hex Addr	7739	30521
x"00",	-- Hex Addr	773A	30522
x"00",	-- Hex Addr	773B	30523
x"00",	-- Hex Addr	773C	30524
x"00",	-- Hex Addr	773D	30525
x"00",	-- Hex Addr	773E	30526
x"00",	-- Hex Addr	773F	30527
x"00",	-- Hex Addr	7740	30528
x"00",	-- Hex Addr	7741	30529
x"00",	-- Hex Addr	7742	30530
x"00",	-- Hex Addr	7743	30531
x"00",	-- Hex Addr	7744	30532
x"00",	-- Hex Addr	7745	30533
x"00",	-- Hex Addr	7746	30534
x"00",	-- Hex Addr	7747	30535
x"00",	-- Hex Addr	7748	30536
x"00",	-- Hex Addr	7749	30537
x"00",	-- Hex Addr	774A	30538
x"00",	-- Hex Addr	774B	30539
x"00",	-- Hex Addr	774C	30540
x"00",	-- Hex Addr	774D	30541
x"00",	-- Hex Addr	774E	30542
x"00",	-- Hex Addr	774F	30543
x"00",	-- Hex Addr	7750	30544
x"00",	-- Hex Addr	7751	30545
x"00",	-- Hex Addr	7752	30546
x"00",	-- Hex Addr	7753	30547
x"00",	-- Hex Addr	7754	30548
x"00",	-- Hex Addr	7755	30549
x"00",	-- Hex Addr	7756	30550
x"00",	-- Hex Addr	7757	30551
x"00",	-- Hex Addr	7758	30552
x"00",	-- Hex Addr	7759	30553
x"00",	-- Hex Addr	775A	30554
x"00",	-- Hex Addr	775B	30555
x"00",	-- Hex Addr	775C	30556
x"00",	-- Hex Addr	775D	30557
x"00",	-- Hex Addr	775E	30558
x"00",	-- Hex Addr	775F	30559
x"00",	-- Hex Addr	7760	30560
x"00",	-- Hex Addr	7761	30561
x"00",	-- Hex Addr	7762	30562
x"00",	-- Hex Addr	7763	30563
x"00",	-- Hex Addr	7764	30564
x"00",	-- Hex Addr	7765	30565
x"00",	-- Hex Addr	7766	30566
x"00",	-- Hex Addr	7767	30567
x"00",	-- Hex Addr	7768	30568
x"00",	-- Hex Addr	7769	30569
x"00",	-- Hex Addr	776A	30570
x"00",	-- Hex Addr	776B	30571
x"00",	-- Hex Addr	776C	30572
x"00",	-- Hex Addr	776D	30573
x"00",	-- Hex Addr	776E	30574
x"00",	-- Hex Addr	776F	30575
x"00",	-- Hex Addr	7770	30576
x"00",	-- Hex Addr	7771	30577
x"00",	-- Hex Addr	7772	30578
x"00",	-- Hex Addr	7773	30579
x"00",	-- Hex Addr	7774	30580
x"00",	-- Hex Addr	7775	30581
x"00",	-- Hex Addr	7776	30582
x"00",	-- Hex Addr	7777	30583
x"00",	-- Hex Addr	7778	30584
x"00",	-- Hex Addr	7779	30585
x"00",	-- Hex Addr	777A	30586
x"00",	-- Hex Addr	777B	30587
x"00",	-- Hex Addr	777C	30588
x"00",	-- Hex Addr	777D	30589
x"00",	-- Hex Addr	777E	30590
x"00",	-- Hex Addr	777F	30591
x"00",	-- Hex Addr	7780	30592
x"00",	-- Hex Addr	7781	30593
x"00",	-- Hex Addr	7782	30594
x"00",	-- Hex Addr	7783	30595
x"00",	-- Hex Addr	7784	30596
x"00",	-- Hex Addr	7785	30597
x"00",	-- Hex Addr	7786	30598
x"00",	-- Hex Addr	7787	30599
x"00",	-- Hex Addr	7788	30600
x"00",	-- Hex Addr	7789	30601
x"00",	-- Hex Addr	778A	30602
x"00",	-- Hex Addr	778B	30603
x"00",	-- Hex Addr	778C	30604
x"00",	-- Hex Addr	778D	30605
x"00",	-- Hex Addr	778E	30606
x"00",	-- Hex Addr	778F	30607
x"00",	-- Hex Addr	7790	30608
x"00",	-- Hex Addr	7791	30609
x"00",	-- Hex Addr	7792	30610
x"00",	-- Hex Addr	7793	30611
x"00",	-- Hex Addr	7794	30612
x"00",	-- Hex Addr	7795	30613
x"00",	-- Hex Addr	7796	30614
x"00",	-- Hex Addr	7797	30615
x"00",	-- Hex Addr	7798	30616
x"00",	-- Hex Addr	7799	30617
x"00",	-- Hex Addr	779A	30618
x"00",	-- Hex Addr	779B	30619
x"00",	-- Hex Addr	779C	30620
x"00",	-- Hex Addr	779D	30621
x"00",	-- Hex Addr	779E	30622
x"00",	-- Hex Addr	779F	30623
x"00",	-- Hex Addr	77A0	30624
x"00",	-- Hex Addr	77A1	30625
x"00",	-- Hex Addr	77A2	30626
x"00",	-- Hex Addr	77A3	30627
x"00",	-- Hex Addr	77A4	30628
x"00",	-- Hex Addr	77A5	30629
x"00",	-- Hex Addr	77A6	30630
x"00",	-- Hex Addr	77A7	30631
x"00",	-- Hex Addr	77A8	30632
x"00",	-- Hex Addr	77A9	30633
x"00",	-- Hex Addr	77AA	30634
x"00",	-- Hex Addr	77AB	30635
x"00",	-- Hex Addr	77AC	30636
x"00",	-- Hex Addr	77AD	30637
x"00",	-- Hex Addr	77AE	30638
x"00",	-- Hex Addr	77AF	30639
x"00",	-- Hex Addr	77B0	30640
x"00",	-- Hex Addr	77B1	30641
x"00",	-- Hex Addr	77B2	30642
x"00",	-- Hex Addr	77B3	30643
x"00",	-- Hex Addr	77B4	30644
x"00",	-- Hex Addr	77B5	30645
x"00",	-- Hex Addr	77B6	30646
x"00",	-- Hex Addr	77B7	30647
x"00",	-- Hex Addr	77B8	30648
x"00",	-- Hex Addr	77B9	30649
x"00",	-- Hex Addr	77BA	30650
x"00",	-- Hex Addr	77BB	30651
x"00",	-- Hex Addr	77BC	30652
x"00",	-- Hex Addr	77BD	30653
x"00",	-- Hex Addr	77BE	30654
x"00",	-- Hex Addr	77BF	30655
x"00",	-- Hex Addr	77C0	30656
x"00",	-- Hex Addr	77C1	30657
x"00",	-- Hex Addr	77C2	30658
x"00",	-- Hex Addr	77C3	30659
x"00",	-- Hex Addr	77C4	30660
x"00",	-- Hex Addr	77C5	30661
x"00",	-- Hex Addr	77C6	30662
x"00",	-- Hex Addr	77C7	30663
x"00",	-- Hex Addr	77C8	30664
x"00",	-- Hex Addr	77C9	30665
x"00",	-- Hex Addr	77CA	30666
x"00",	-- Hex Addr	77CB	30667
x"00",	-- Hex Addr	77CC	30668
x"00",	-- Hex Addr	77CD	30669
x"00",	-- Hex Addr	77CE	30670
x"00",	-- Hex Addr	77CF	30671
x"00",	-- Hex Addr	77D0	30672
x"00",	-- Hex Addr	77D1	30673
x"00",	-- Hex Addr	77D2	30674
x"00",	-- Hex Addr	77D3	30675
x"00",	-- Hex Addr	77D4	30676
x"00",	-- Hex Addr	77D5	30677
x"00",	-- Hex Addr	77D6	30678
x"00",	-- Hex Addr	77D7	30679
x"00",	-- Hex Addr	77D8	30680
x"00",	-- Hex Addr	77D9	30681
x"00",	-- Hex Addr	77DA	30682
x"00",	-- Hex Addr	77DB	30683
x"00",	-- Hex Addr	77DC	30684
x"00",	-- Hex Addr	77DD	30685
x"00",	-- Hex Addr	77DE	30686
x"00",	-- Hex Addr	77DF	30687
x"00",	-- Hex Addr	77E0	30688
x"00",	-- Hex Addr	77E1	30689
x"00",	-- Hex Addr	77E2	30690
x"00",	-- Hex Addr	77E3	30691
x"00",	-- Hex Addr	77E4	30692
x"00",	-- Hex Addr	77E5	30693
x"00",	-- Hex Addr	77E6	30694
x"00",	-- Hex Addr	77E7	30695
x"00",	-- Hex Addr	77E8	30696
x"00",	-- Hex Addr	77E9	30697
x"00",	-- Hex Addr	77EA	30698
x"00",	-- Hex Addr	77EB	30699
x"00",	-- Hex Addr	77EC	30700
x"00",	-- Hex Addr	77ED	30701
x"00",	-- Hex Addr	77EE	30702
x"00",	-- Hex Addr	77EF	30703
x"00",	-- Hex Addr	77F0	30704
x"00",	-- Hex Addr	77F1	30705
x"00",	-- Hex Addr	77F2	30706
x"00",	-- Hex Addr	77F3	30707
x"00",	-- Hex Addr	77F4	30708
x"00",	-- Hex Addr	77F5	30709
x"00",	-- Hex Addr	77F6	30710
x"00",	-- Hex Addr	77F7	30711
x"00",	-- Hex Addr	77F8	30712
x"00",	-- Hex Addr	77F9	30713
x"00",	-- Hex Addr	77FA	30714
x"00",	-- Hex Addr	77FB	30715
x"00",	-- Hex Addr	77FC	30716
x"00",	-- Hex Addr	77FD	30717
x"00",	-- Hex Addr	77FE	30718
x"00",	-- Hex Addr	77FF	30719
x"00",	-- Hex Addr	7800	30720
x"00",	-- Hex Addr	7801	30721
x"00",	-- Hex Addr	7802	30722
x"00",	-- Hex Addr	7803	30723
x"00",	-- Hex Addr	7804	30724
x"00",	-- Hex Addr	7805	30725
x"00",	-- Hex Addr	7806	30726
x"00",	-- Hex Addr	7807	30727
x"00",	-- Hex Addr	7808	30728
x"00",	-- Hex Addr	7809	30729
x"00",	-- Hex Addr	780A	30730
x"00",	-- Hex Addr	780B	30731
x"00",	-- Hex Addr	780C	30732
x"00",	-- Hex Addr	780D	30733
x"00",	-- Hex Addr	780E	30734
x"00",	-- Hex Addr	780F	30735
x"00",	-- Hex Addr	7810	30736
x"00",	-- Hex Addr	7811	30737
x"00",	-- Hex Addr	7812	30738
x"00",	-- Hex Addr	7813	30739
x"00",	-- Hex Addr	7814	30740
x"00",	-- Hex Addr	7815	30741
x"00",	-- Hex Addr	7816	30742
x"00",	-- Hex Addr	7817	30743
x"00",	-- Hex Addr	7818	30744
x"00",	-- Hex Addr	7819	30745
x"00",	-- Hex Addr	781A	30746
x"00",	-- Hex Addr	781B	30747
x"00",	-- Hex Addr	781C	30748
x"00",	-- Hex Addr	781D	30749
x"00",	-- Hex Addr	781E	30750
x"00",	-- Hex Addr	781F	30751
x"00",	-- Hex Addr	7820	30752
x"00",	-- Hex Addr	7821	30753
x"00",	-- Hex Addr	7822	30754
x"00",	-- Hex Addr	7823	30755
x"00",	-- Hex Addr	7824	30756
x"00",	-- Hex Addr	7825	30757
x"00",	-- Hex Addr	7826	30758
x"00",	-- Hex Addr	7827	30759
x"00",	-- Hex Addr	7828	30760
x"00",	-- Hex Addr	7829	30761
x"00",	-- Hex Addr	782A	30762
x"00",	-- Hex Addr	782B	30763
x"00",	-- Hex Addr	782C	30764
x"00",	-- Hex Addr	782D	30765
x"00",	-- Hex Addr	782E	30766
x"00",	-- Hex Addr	782F	30767
x"00",	-- Hex Addr	7830	30768
x"00",	-- Hex Addr	7831	30769
x"00",	-- Hex Addr	7832	30770
x"00",	-- Hex Addr	7833	30771
x"00",	-- Hex Addr	7834	30772
x"00",	-- Hex Addr	7835	30773
x"00",	-- Hex Addr	7836	30774
x"00",	-- Hex Addr	7837	30775
x"00",	-- Hex Addr	7838	30776
x"00",	-- Hex Addr	7839	30777
x"00",	-- Hex Addr	783A	30778
x"00",	-- Hex Addr	783B	30779
x"00",	-- Hex Addr	783C	30780
x"00",	-- Hex Addr	783D	30781
x"00",	-- Hex Addr	783E	30782
x"00",	-- Hex Addr	783F	30783
x"00",	-- Hex Addr	7840	30784
x"00",	-- Hex Addr	7841	30785
x"00",	-- Hex Addr	7842	30786
x"00",	-- Hex Addr	7843	30787
x"00",	-- Hex Addr	7844	30788
x"00",	-- Hex Addr	7845	30789
x"00",	-- Hex Addr	7846	30790
x"00",	-- Hex Addr	7847	30791
x"00",	-- Hex Addr	7848	30792
x"00",	-- Hex Addr	7849	30793
x"00",	-- Hex Addr	784A	30794
x"00",	-- Hex Addr	784B	30795
x"00",	-- Hex Addr	784C	30796
x"00",	-- Hex Addr	784D	30797
x"00",	-- Hex Addr	784E	30798
x"00",	-- Hex Addr	784F	30799
x"00",	-- Hex Addr	7850	30800
x"00",	-- Hex Addr	7851	30801
x"00",	-- Hex Addr	7852	30802
x"00",	-- Hex Addr	7853	30803
x"00",	-- Hex Addr	7854	30804
x"00",	-- Hex Addr	7855	30805
x"00",	-- Hex Addr	7856	30806
x"00",	-- Hex Addr	7857	30807
x"00",	-- Hex Addr	7858	30808
x"00",	-- Hex Addr	7859	30809
x"00",	-- Hex Addr	785A	30810
x"00",	-- Hex Addr	785B	30811
x"00",	-- Hex Addr	785C	30812
x"00",	-- Hex Addr	785D	30813
x"00",	-- Hex Addr	785E	30814
x"00",	-- Hex Addr	785F	30815
x"00",	-- Hex Addr	7860	30816
x"00",	-- Hex Addr	7861	30817
x"00",	-- Hex Addr	7862	30818
x"00",	-- Hex Addr	7863	30819
x"00",	-- Hex Addr	7864	30820
x"00",	-- Hex Addr	7865	30821
x"00",	-- Hex Addr	7866	30822
x"00",	-- Hex Addr	7867	30823
x"00",	-- Hex Addr	7868	30824
x"00",	-- Hex Addr	7869	30825
x"00",	-- Hex Addr	786A	30826
x"00",	-- Hex Addr	786B	30827
x"00",	-- Hex Addr	786C	30828
x"00",	-- Hex Addr	786D	30829
x"00",	-- Hex Addr	786E	30830
x"00",	-- Hex Addr	786F	30831
x"00",	-- Hex Addr	7870	30832
x"00",	-- Hex Addr	7871	30833
x"00",	-- Hex Addr	7872	30834
x"00",	-- Hex Addr	7873	30835
x"00",	-- Hex Addr	7874	30836
x"00",	-- Hex Addr	7875	30837
x"00",	-- Hex Addr	7876	30838
x"00",	-- Hex Addr	7877	30839
x"00",	-- Hex Addr	7878	30840
x"00",	-- Hex Addr	7879	30841
x"00",	-- Hex Addr	787A	30842
x"00",	-- Hex Addr	787B	30843
x"00",	-- Hex Addr	787C	30844
x"00",	-- Hex Addr	787D	30845
x"00",	-- Hex Addr	787E	30846
x"00",	-- Hex Addr	787F	30847
x"00",	-- Hex Addr	7880	30848
x"00",	-- Hex Addr	7881	30849
x"00",	-- Hex Addr	7882	30850
x"00",	-- Hex Addr	7883	30851
x"00",	-- Hex Addr	7884	30852
x"00",	-- Hex Addr	7885	30853
x"00",	-- Hex Addr	7886	30854
x"00",	-- Hex Addr	7887	30855
x"00",	-- Hex Addr	7888	30856
x"00",	-- Hex Addr	7889	30857
x"00",	-- Hex Addr	788A	30858
x"00",	-- Hex Addr	788B	30859
x"00",	-- Hex Addr	788C	30860
x"00",	-- Hex Addr	788D	30861
x"00",	-- Hex Addr	788E	30862
x"00",	-- Hex Addr	788F	30863
x"00",	-- Hex Addr	7890	30864
x"00",	-- Hex Addr	7891	30865
x"00",	-- Hex Addr	7892	30866
x"00",	-- Hex Addr	7893	30867
x"00",	-- Hex Addr	7894	30868
x"00",	-- Hex Addr	7895	30869
x"00",	-- Hex Addr	7896	30870
x"00",	-- Hex Addr	7897	30871
x"00",	-- Hex Addr	7898	30872
x"00",	-- Hex Addr	7899	30873
x"00",	-- Hex Addr	789A	30874
x"00",	-- Hex Addr	789B	30875
x"00",	-- Hex Addr	789C	30876
x"00",	-- Hex Addr	789D	30877
x"00",	-- Hex Addr	789E	30878
x"00",	-- Hex Addr	789F	30879
x"00",	-- Hex Addr	78A0	30880
x"00",	-- Hex Addr	78A1	30881
x"00",	-- Hex Addr	78A2	30882
x"00",	-- Hex Addr	78A3	30883
x"00",	-- Hex Addr	78A4	30884
x"00",	-- Hex Addr	78A5	30885
x"00",	-- Hex Addr	78A6	30886
x"00",	-- Hex Addr	78A7	30887
x"00",	-- Hex Addr	78A8	30888
x"00",	-- Hex Addr	78A9	30889
x"00",	-- Hex Addr	78AA	30890
x"00",	-- Hex Addr	78AB	30891
x"00",	-- Hex Addr	78AC	30892
x"00",	-- Hex Addr	78AD	30893
x"00",	-- Hex Addr	78AE	30894
x"00",	-- Hex Addr	78AF	30895
x"00",	-- Hex Addr	78B0	30896
x"00",	-- Hex Addr	78B1	30897
x"00",	-- Hex Addr	78B2	30898
x"00",	-- Hex Addr	78B3	30899
x"00",	-- Hex Addr	78B4	30900
x"00",	-- Hex Addr	78B5	30901
x"00",	-- Hex Addr	78B6	30902
x"00",	-- Hex Addr	78B7	30903
x"00",	-- Hex Addr	78B8	30904
x"00",	-- Hex Addr	78B9	30905
x"00",	-- Hex Addr	78BA	30906
x"00",	-- Hex Addr	78BB	30907
x"00",	-- Hex Addr	78BC	30908
x"00",	-- Hex Addr	78BD	30909
x"00",	-- Hex Addr	78BE	30910
x"00",	-- Hex Addr	78BF	30911
x"00",	-- Hex Addr	78C0	30912
x"00",	-- Hex Addr	78C1	30913
x"00",	-- Hex Addr	78C2	30914
x"00",	-- Hex Addr	78C3	30915
x"00",	-- Hex Addr	78C4	30916
x"00",	-- Hex Addr	78C5	30917
x"00",	-- Hex Addr	78C6	30918
x"00",	-- Hex Addr	78C7	30919
x"00",	-- Hex Addr	78C8	30920
x"00",	-- Hex Addr	78C9	30921
x"00",	-- Hex Addr	78CA	30922
x"00",	-- Hex Addr	78CB	30923
x"00",	-- Hex Addr	78CC	30924
x"00",	-- Hex Addr	78CD	30925
x"00",	-- Hex Addr	78CE	30926
x"00",	-- Hex Addr	78CF	30927
x"00",	-- Hex Addr	78D0	30928
x"00",	-- Hex Addr	78D1	30929
x"00",	-- Hex Addr	78D2	30930
x"00",	-- Hex Addr	78D3	30931
x"00",	-- Hex Addr	78D4	30932
x"00",	-- Hex Addr	78D5	30933
x"00",	-- Hex Addr	78D6	30934
x"00",	-- Hex Addr	78D7	30935
x"00",	-- Hex Addr	78D8	30936
x"00",	-- Hex Addr	78D9	30937
x"00",	-- Hex Addr	78DA	30938
x"00",	-- Hex Addr	78DB	30939
x"00",	-- Hex Addr	78DC	30940
x"00",	-- Hex Addr	78DD	30941
x"00",	-- Hex Addr	78DE	30942
x"00",	-- Hex Addr	78DF	30943
x"00",	-- Hex Addr	78E0	30944
x"00",	-- Hex Addr	78E1	30945
x"00",	-- Hex Addr	78E2	30946
x"00",	-- Hex Addr	78E3	30947
x"00",	-- Hex Addr	78E4	30948
x"00",	-- Hex Addr	78E5	30949
x"00",	-- Hex Addr	78E6	30950
x"00",	-- Hex Addr	78E7	30951
x"00",	-- Hex Addr	78E8	30952
x"00",	-- Hex Addr	78E9	30953
x"00",	-- Hex Addr	78EA	30954
x"00",	-- Hex Addr	78EB	30955
x"00",	-- Hex Addr	78EC	30956
x"00",	-- Hex Addr	78ED	30957
x"00",	-- Hex Addr	78EE	30958
x"00",	-- Hex Addr	78EF	30959
x"00",	-- Hex Addr	78F0	30960
x"00",	-- Hex Addr	78F1	30961
x"00",	-- Hex Addr	78F2	30962
x"00",	-- Hex Addr	78F3	30963
x"00",	-- Hex Addr	78F4	30964
x"00",	-- Hex Addr	78F5	30965
x"00",	-- Hex Addr	78F6	30966
x"00",	-- Hex Addr	78F7	30967
x"00",	-- Hex Addr	78F8	30968
x"00",	-- Hex Addr	78F9	30969
x"00",	-- Hex Addr	78FA	30970
x"00",	-- Hex Addr	78FB	30971
x"00",	-- Hex Addr	78FC	30972
x"00",	-- Hex Addr	78FD	30973
x"00",	-- Hex Addr	78FE	30974
x"00",	-- Hex Addr	78FF	30975
x"00",	-- Hex Addr	7900	30976
x"00",	-- Hex Addr	7901	30977
x"00",	-- Hex Addr	7902	30978
x"00",	-- Hex Addr	7903	30979
x"00",	-- Hex Addr	7904	30980
x"00",	-- Hex Addr	7905	30981
x"00",	-- Hex Addr	7906	30982
x"00",	-- Hex Addr	7907	30983
x"00",	-- Hex Addr	7908	30984
x"00",	-- Hex Addr	7909	30985
x"00",	-- Hex Addr	790A	30986
x"00",	-- Hex Addr	790B	30987
x"00",	-- Hex Addr	790C	30988
x"00",	-- Hex Addr	790D	30989
x"00",	-- Hex Addr	790E	30990
x"00",	-- Hex Addr	790F	30991
x"00",	-- Hex Addr	7910	30992
x"00",	-- Hex Addr	7911	30993
x"00",	-- Hex Addr	7912	30994
x"00",	-- Hex Addr	7913	30995
x"00",	-- Hex Addr	7914	30996
x"00",	-- Hex Addr	7915	30997
x"00",	-- Hex Addr	7916	30998
x"00",	-- Hex Addr	7917	30999
x"00",	-- Hex Addr	7918	31000
x"00",	-- Hex Addr	7919	31001
x"00",	-- Hex Addr	791A	31002
x"00",	-- Hex Addr	791B	31003
x"00",	-- Hex Addr	791C	31004
x"00",	-- Hex Addr	791D	31005
x"00",	-- Hex Addr	791E	31006
x"00",	-- Hex Addr	791F	31007
x"00",	-- Hex Addr	7920	31008
x"00",	-- Hex Addr	7921	31009
x"00",	-- Hex Addr	7922	31010
x"00",	-- Hex Addr	7923	31011
x"00",	-- Hex Addr	7924	31012
x"00",	-- Hex Addr	7925	31013
x"00",	-- Hex Addr	7926	31014
x"00",	-- Hex Addr	7927	31015
x"00",	-- Hex Addr	7928	31016
x"00",	-- Hex Addr	7929	31017
x"00",	-- Hex Addr	792A	31018
x"00",	-- Hex Addr	792B	31019
x"00",	-- Hex Addr	792C	31020
x"00",	-- Hex Addr	792D	31021
x"00",	-- Hex Addr	792E	31022
x"00",	-- Hex Addr	792F	31023
x"00",	-- Hex Addr	7930	31024
x"00",	-- Hex Addr	7931	31025
x"00",	-- Hex Addr	7932	31026
x"00",	-- Hex Addr	7933	31027
x"00",	-- Hex Addr	7934	31028
x"00",	-- Hex Addr	7935	31029
x"00",	-- Hex Addr	7936	31030
x"00",	-- Hex Addr	7937	31031
x"00",	-- Hex Addr	7938	31032
x"00",	-- Hex Addr	7939	31033
x"00",	-- Hex Addr	793A	31034
x"00",	-- Hex Addr	793B	31035
x"00",	-- Hex Addr	793C	31036
x"00",	-- Hex Addr	793D	31037
x"00",	-- Hex Addr	793E	31038
x"00",	-- Hex Addr	793F	31039
x"00",	-- Hex Addr	7940	31040
x"00",	-- Hex Addr	7941	31041
x"00",	-- Hex Addr	7942	31042
x"00",	-- Hex Addr	7943	31043
x"00",	-- Hex Addr	7944	31044
x"00",	-- Hex Addr	7945	31045
x"00",	-- Hex Addr	7946	31046
x"00",	-- Hex Addr	7947	31047
x"00",	-- Hex Addr	7948	31048
x"00",	-- Hex Addr	7949	31049
x"00",	-- Hex Addr	794A	31050
x"00",	-- Hex Addr	794B	31051
x"00",	-- Hex Addr	794C	31052
x"00",	-- Hex Addr	794D	31053
x"00",	-- Hex Addr	794E	31054
x"00",	-- Hex Addr	794F	31055
x"00",	-- Hex Addr	7950	31056
x"00",	-- Hex Addr	7951	31057
x"00",	-- Hex Addr	7952	31058
x"00",	-- Hex Addr	7953	31059
x"00",	-- Hex Addr	7954	31060
x"00",	-- Hex Addr	7955	31061
x"00",	-- Hex Addr	7956	31062
x"00",	-- Hex Addr	7957	31063
x"00",	-- Hex Addr	7958	31064
x"00",	-- Hex Addr	7959	31065
x"00",	-- Hex Addr	795A	31066
x"00",	-- Hex Addr	795B	31067
x"00",	-- Hex Addr	795C	31068
x"00",	-- Hex Addr	795D	31069
x"00",	-- Hex Addr	795E	31070
x"00",	-- Hex Addr	795F	31071
x"00",	-- Hex Addr	7960	31072
x"00",	-- Hex Addr	7961	31073
x"00",	-- Hex Addr	7962	31074
x"00",	-- Hex Addr	7963	31075
x"00",	-- Hex Addr	7964	31076
x"00",	-- Hex Addr	7965	31077
x"00",	-- Hex Addr	7966	31078
x"00",	-- Hex Addr	7967	31079
x"00",	-- Hex Addr	7968	31080
x"00",	-- Hex Addr	7969	31081
x"00",	-- Hex Addr	796A	31082
x"00",	-- Hex Addr	796B	31083
x"00",	-- Hex Addr	796C	31084
x"00",	-- Hex Addr	796D	31085
x"00",	-- Hex Addr	796E	31086
x"00",	-- Hex Addr	796F	31087
x"00",	-- Hex Addr	7970	31088
x"00",	-- Hex Addr	7971	31089
x"00",	-- Hex Addr	7972	31090
x"00",	-- Hex Addr	7973	31091
x"00",	-- Hex Addr	7974	31092
x"00",	-- Hex Addr	7975	31093
x"00",	-- Hex Addr	7976	31094
x"00",	-- Hex Addr	7977	31095
x"00",	-- Hex Addr	7978	31096
x"00",	-- Hex Addr	7979	31097
x"00",	-- Hex Addr	797A	31098
x"00",	-- Hex Addr	797B	31099
x"00",	-- Hex Addr	797C	31100
x"00",	-- Hex Addr	797D	31101
x"00",	-- Hex Addr	797E	31102
x"00",	-- Hex Addr	797F	31103
x"00",	-- Hex Addr	7980	31104
x"00",	-- Hex Addr	7981	31105
x"00",	-- Hex Addr	7982	31106
x"00",	-- Hex Addr	7983	31107
x"00",	-- Hex Addr	7984	31108
x"00",	-- Hex Addr	7985	31109
x"00",	-- Hex Addr	7986	31110
x"00",	-- Hex Addr	7987	31111
x"00",	-- Hex Addr	7988	31112
x"00",	-- Hex Addr	7989	31113
x"00",	-- Hex Addr	798A	31114
x"00",	-- Hex Addr	798B	31115
x"00",	-- Hex Addr	798C	31116
x"00",	-- Hex Addr	798D	31117
x"00",	-- Hex Addr	798E	31118
x"00",	-- Hex Addr	798F	31119
x"00",	-- Hex Addr	7990	31120
x"00",	-- Hex Addr	7991	31121
x"00",	-- Hex Addr	7992	31122
x"00",	-- Hex Addr	7993	31123
x"00",	-- Hex Addr	7994	31124
x"00",	-- Hex Addr	7995	31125
x"00",	-- Hex Addr	7996	31126
x"00",	-- Hex Addr	7997	31127
x"00",	-- Hex Addr	7998	31128
x"00",	-- Hex Addr	7999	31129
x"00",	-- Hex Addr	799A	31130
x"00",	-- Hex Addr	799B	31131
x"00",	-- Hex Addr	799C	31132
x"00",	-- Hex Addr	799D	31133
x"00",	-- Hex Addr	799E	31134
x"00",	-- Hex Addr	799F	31135
x"00",	-- Hex Addr	79A0	31136
x"00",	-- Hex Addr	79A1	31137
x"00",	-- Hex Addr	79A2	31138
x"00",	-- Hex Addr	79A3	31139
x"00",	-- Hex Addr	79A4	31140
x"00",	-- Hex Addr	79A5	31141
x"00",	-- Hex Addr	79A6	31142
x"00",	-- Hex Addr	79A7	31143
x"00",	-- Hex Addr	79A8	31144
x"00",	-- Hex Addr	79A9	31145
x"00",	-- Hex Addr	79AA	31146
x"00",	-- Hex Addr	79AB	31147
x"00",	-- Hex Addr	79AC	31148
x"00",	-- Hex Addr	79AD	31149
x"00",	-- Hex Addr	79AE	31150
x"00",	-- Hex Addr	79AF	31151
x"00",	-- Hex Addr	79B0	31152
x"00",	-- Hex Addr	79B1	31153
x"00",	-- Hex Addr	79B2	31154
x"00",	-- Hex Addr	79B3	31155
x"00",	-- Hex Addr	79B4	31156
x"00",	-- Hex Addr	79B5	31157
x"00",	-- Hex Addr	79B6	31158
x"00",	-- Hex Addr	79B7	31159
x"00",	-- Hex Addr	79B8	31160
x"00",	-- Hex Addr	79B9	31161
x"00",	-- Hex Addr	79BA	31162
x"00",	-- Hex Addr	79BB	31163
x"00",	-- Hex Addr	79BC	31164
x"00",	-- Hex Addr	79BD	31165
x"00",	-- Hex Addr	79BE	31166
x"00",	-- Hex Addr	79BF	31167
x"00",	-- Hex Addr	79C0	31168
x"00",	-- Hex Addr	79C1	31169
x"00",	-- Hex Addr	79C2	31170
x"00",	-- Hex Addr	79C3	31171
x"00",	-- Hex Addr	79C4	31172
x"00",	-- Hex Addr	79C5	31173
x"00",	-- Hex Addr	79C6	31174
x"00",	-- Hex Addr	79C7	31175
x"00",	-- Hex Addr	79C8	31176
x"00",	-- Hex Addr	79C9	31177
x"00",	-- Hex Addr	79CA	31178
x"00",	-- Hex Addr	79CB	31179
x"00",	-- Hex Addr	79CC	31180
x"00",	-- Hex Addr	79CD	31181
x"00",	-- Hex Addr	79CE	31182
x"00",	-- Hex Addr	79CF	31183
x"00",	-- Hex Addr	79D0	31184
x"00",	-- Hex Addr	79D1	31185
x"00",	-- Hex Addr	79D2	31186
x"00",	-- Hex Addr	79D3	31187
x"00",	-- Hex Addr	79D4	31188
x"00",	-- Hex Addr	79D5	31189
x"00",	-- Hex Addr	79D6	31190
x"00",	-- Hex Addr	79D7	31191
x"00",	-- Hex Addr	79D8	31192
x"00",	-- Hex Addr	79D9	31193
x"00",	-- Hex Addr	79DA	31194
x"00",	-- Hex Addr	79DB	31195
x"00",	-- Hex Addr	79DC	31196
x"00",	-- Hex Addr	79DD	31197
x"00",	-- Hex Addr	79DE	31198
x"00",	-- Hex Addr	79DF	31199
x"00",	-- Hex Addr	79E0	31200
x"00",	-- Hex Addr	79E1	31201
x"00",	-- Hex Addr	79E2	31202
x"00",	-- Hex Addr	79E3	31203
x"00",	-- Hex Addr	79E4	31204
x"00",	-- Hex Addr	79E5	31205
x"00",	-- Hex Addr	79E6	31206
x"00",	-- Hex Addr	79E7	31207
x"00",	-- Hex Addr	79E8	31208
x"00",	-- Hex Addr	79E9	31209
x"00",	-- Hex Addr	79EA	31210
x"00",	-- Hex Addr	79EB	31211
x"00",	-- Hex Addr	79EC	31212
x"00",	-- Hex Addr	79ED	31213
x"00",	-- Hex Addr	79EE	31214
x"00",	-- Hex Addr	79EF	31215
x"00",	-- Hex Addr	79F0	31216
x"00",	-- Hex Addr	79F1	31217
x"00",	-- Hex Addr	79F2	31218
x"00",	-- Hex Addr	79F3	31219
x"00",	-- Hex Addr	79F4	31220
x"00",	-- Hex Addr	79F5	31221
x"00",	-- Hex Addr	79F6	31222
x"00",	-- Hex Addr	79F7	31223
x"00",	-- Hex Addr	79F8	31224
x"00",	-- Hex Addr	79F9	31225
x"00",	-- Hex Addr	79FA	31226
x"00",	-- Hex Addr	79FB	31227
x"00",	-- Hex Addr	79FC	31228
x"00",	-- Hex Addr	79FD	31229
x"00",	-- Hex Addr	79FE	31230
x"00",	-- Hex Addr	79FF	31231
x"00",	-- Hex Addr	7A00	31232
x"00",	-- Hex Addr	7A01	31233
x"00",	-- Hex Addr	7A02	31234
x"00",	-- Hex Addr	7A03	31235
x"00",	-- Hex Addr	7A04	31236
x"00",	-- Hex Addr	7A05	31237
x"00",	-- Hex Addr	7A06	31238
x"00",	-- Hex Addr	7A07	31239
x"00",	-- Hex Addr	7A08	31240
x"00",	-- Hex Addr	7A09	31241
x"00",	-- Hex Addr	7A0A	31242
x"00",	-- Hex Addr	7A0B	31243
x"00",	-- Hex Addr	7A0C	31244
x"00",	-- Hex Addr	7A0D	31245
x"00",	-- Hex Addr	7A0E	31246
x"00",	-- Hex Addr	7A0F	31247
x"00",	-- Hex Addr	7A10	31248
x"00",	-- Hex Addr	7A11	31249
x"00",	-- Hex Addr	7A12	31250
x"00",	-- Hex Addr	7A13	31251
x"00",	-- Hex Addr	7A14	31252
x"00",	-- Hex Addr	7A15	31253
x"00",	-- Hex Addr	7A16	31254
x"00",	-- Hex Addr	7A17	31255
x"00",	-- Hex Addr	7A18	31256
x"00",	-- Hex Addr	7A19	31257
x"00",	-- Hex Addr	7A1A	31258
x"00",	-- Hex Addr	7A1B	31259
x"00",	-- Hex Addr	7A1C	31260
x"00",	-- Hex Addr	7A1D	31261
x"00",	-- Hex Addr	7A1E	31262
x"00",	-- Hex Addr	7A1F	31263
x"00",	-- Hex Addr	7A20	31264
x"00",	-- Hex Addr	7A21	31265
x"00",	-- Hex Addr	7A22	31266
x"00",	-- Hex Addr	7A23	31267
x"00",	-- Hex Addr	7A24	31268
x"00",	-- Hex Addr	7A25	31269
x"00",	-- Hex Addr	7A26	31270
x"00",	-- Hex Addr	7A27	31271
x"00",	-- Hex Addr	7A28	31272
x"00",	-- Hex Addr	7A29	31273
x"00",	-- Hex Addr	7A2A	31274
x"00",	-- Hex Addr	7A2B	31275
x"00",	-- Hex Addr	7A2C	31276
x"00",	-- Hex Addr	7A2D	31277
x"00",	-- Hex Addr	7A2E	31278
x"00",	-- Hex Addr	7A2F	31279
x"00",	-- Hex Addr	7A30	31280
x"00",	-- Hex Addr	7A31	31281
x"00",	-- Hex Addr	7A32	31282
x"00",	-- Hex Addr	7A33	31283
x"00",	-- Hex Addr	7A34	31284
x"00",	-- Hex Addr	7A35	31285
x"00",	-- Hex Addr	7A36	31286
x"00",	-- Hex Addr	7A37	31287
x"00",	-- Hex Addr	7A38	31288
x"00",	-- Hex Addr	7A39	31289
x"00",	-- Hex Addr	7A3A	31290
x"00",	-- Hex Addr	7A3B	31291
x"00",	-- Hex Addr	7A3C	31292
x"00",	-- Hex Addr	7A3D	31293
x"00",	-- Hex Addr	7A3E	31294
x"00",	-- Hex Addr	7A3F	31295
x"00",	-- Hex Addr	7A40	31296
x"00",	-- Hex Addr	7A41	31297
x"00",	-- Hex Addr	7A42	31298
x"00",	-- Hex Addr	7A43	31299
x"00",	-- Hex Addr	7A44	31300
x"00",	-- Hex Addr	7A45	31301
x"00",	-- Hex Addr	7A46	31302
x"00",	-- Hex Addr	7A47	31303
x"00",	-- Hex Addr	7A48	31304
x"00",	-- Hex Addr	7A49	31305
x"00",	-- Hex Addr	7A4A	31306
x"00",	-- Hex Addr	7A4B	31307
x"00",	-- Hex Addr	7A4C	31308
x"00",	-- Hex Addr	7A4D	31309
x"00",	-- Hex Addr	7A4E	31310
x"00",	-- Hex Addr	7A4F	31311
x"00",	-- Hex Addr	7A50	31312
x"00",	-- Hex Addr	7A51	31313
x"00",	-- Hex Addr	7A52	31314
x"00",	-- Hex Addr	7A53	31315
x"00",	-- Hex Addr	7A54	31316
x"00",	-- Hex Addr	7A55	31317
x"00",	-- Hex Addr	7A56	31318
x"00",	-- Hex Addr	7A57	31319
x"00",	-- Hex Addr	7A58	31320
x"00",	-- Hex Addr	7A59	31321
x"00",	-- Hex Addr	7A5A	31322
x"00",	-- Hex Addr	7A5B	31323
x"00",	-- Hex Addr	7A5C	31324
x"00",	-- Hex Addr	7A5D	31325
x"00",	-- Hex Addr	7A5E	31326
x"00",	-- Hex Addr	7A5F	31327
x"00",	-- Hex Addr	7A60	31328
x"00",	-- Hex Addr	7A61	31329
x"00",	-- Hex Addr	7A62	31330
x"00",	-- Hex Addr	7A63	31331
x"00",	-- Hex Addr	7A64	31332
x"00",	-- Hex Addr	7A65	31333
x"00",	-- Hex Addr	7A66	31334
x"00",	-- Hex Addr	7A67	31335
x"00",	-- Hex Addr	7A68	31336
x"00",	-- Hex Addr	7A69	31337
x"00",	-- Hex Addr	7A6A	31338
x"00",	-- Hex Addr	7A6B	31339
x"00",	-- Hex Addr	7A6C	31340
x"00",	-- Hex Addr	7A6D	31341
x"00",	-- Hex Addr	7A6E	31342
x"00",	-- Hex Addr	7A6F	31343
x"00",	-- Hex Addr	7A70	31344
x"00",	-- Hex Addr	7A71	31345
x"00",	-- Hex Addr	7A72	31346
x"00",	-- Hex Addr	7A73	31347
x"00",	-- Hex Addr	7A74	31348
x"00",	-- Hex Addr	7A75	31349
x"00",	-- Hex Addr	7A76	31350
x"00",	-- Hex Addr	7A77	31351
x"00",	-- Hex Addr	7A78	31352
x"00",	-- Hex Addr	7A79	31353
x"00",	-- Hex Addr	7A7A	31354
x"00",	-- Hex Addr	7A7B	31355
x"00",	-- Hex Addr	7A7C	31356
x"00",	-- Hex Addr	7A7D	31357
x"00",	-- Hex Addr	7A7E	31358
x"00",	-- Hex Addr	7A7F	31359
x"00",	-- Hex Addr	7A80	31360
x"00",	-- Hex Addr	7A81	31361
x"00",	-- Hex Addr	7A82	31362
x"00",	-- Hex Addr	7A83	31363
x"00",	-- Hex Addr	7A84	31364
x"00",	-- Hex Addr	7A85	31365
x"00",	-- Hex Addr	7A86	31366
x"00",	-- Hex Addr	7A87	31367
x"00",	-- Hex Addr	7A88	31368
x"00",	-- Hex Addr	7A89	31369
x"00",	-- Hex Addr	7A8A	31370
x"00",	-- Hex Addr	7A8B	31371
x"00",	-- Hex Addr	7A8C	31372
x"00",	-- Hex Addr	7A8D	31373
x"00",	-- Hex Addr	7A8E	31374
x"00",	-- Hex Addr	7A8F	31375
x"00",	-- Hex Addr	7A90	31376
x"00",	-- Hex Addr	7A91	31377
x"00",	-- Hex Addr	7A92	31378
x"00",	-- Hex Addr	7A93	31379
x"00",	-- Hex Addr	7A94	31380
x"00",	-- Hex Addr	7A95	31381
x"00",	-- Hex Addr	7A96	31382
x"00",	-- Hex Addr	7A97	31383
x"00",	-- Hex Addr	7A98	31384
x"00",	-- Hex Addr	7A99	31385
x"00",	-- Hex Addr	7A9A	31386
x"00",	-- Hex Addr	7A9B	31387
x"00",	-- Hex Addr	7A9C	31388
x"00",	-- Hex Addr	7A9D	31389
x"00",	-- Hex Addr	7A9E	31390
x"00",	-- Hex Addr	7A9F	31391
x"00",	-- Hex Addr	7AA0	31392
x"00",	-- Hex Addr	7AA1	31393
x"00",	-- Hex Addr	7AA2	31394
x"00",	-- Hex Addr	7AA3	31395
x"00",	-- Hex Addr	7AA4	31396
x"00",	-- Hex Addr	7AA5	31397
x"00",	-- Hex Addr	7AA6	31398
x"00",	-- Hex Addr	7AA7	31399
x"00",	-- Hex Addr	7AA8	31400
x"00",	-- Hex Addr	7AA9	31401
x"00",	-- Hex Addr	7AAA	31402
x"00",	-- Hex Addr	7AAB	31403
x"00",	-- Hex Addr	7AAC	31404
x"00",	-- Hex Addr	7AAD	31405
x"00",	-- Hex Addr	7AAE	31406
x"00",	-- Hex Addr	7AAF	31407
x"00",	-- Hex Addr	7AB0	31408
x"00",	-- Hex Addr	7AB1	31409
x"00",	-- Hex Addr	7AB2	31410
x"00",	-- Hex Addr	7AB3	31411
x"00",	-- Hex Addr	7AB4	31412
x"00",	-- Hex Addr	7AB5	31413
x"00",	-- Hex Addr	7AB6	31414
x"00",	-- Hex Addr	7AB7	31415
x"00",	-- Hex Addr	7AB8	31416
x"00",	-- Hex Addr	7AB9	31417
x"00",	-- Hex Addr	7ABA	31418
x"00",	-- Hex Addr	7ABB	31419
x"00",	-- Hex Addr	7ABC	31420
x"00",	-- Hex Addr	7ABD	31421
x"00",	-- Hex Addr	7ABE	31422
x"00",	-- Hex Addr	7ABF	31423
x"00",	-- Hex Addr	7AC0	31424
x"00",	-- Hex Addr	7AC1	31425
x"00",	-- Hex Addr	7AC2	31426
x"00",	-- Hex Addr	7AC3	31427
x"00",	-- Hex Addr	7AC4	31428
x"00",	-- Hex Addr	7AC5	31429
x"00",	-- Hex Addr	7AC6	31430
x"00",	-- Hex Addr	7AC7	31431
x"00",	-- Hex Addr	7AC8	31432
x"00",	-- Hex Addr	7AC9	31433
x"00",	-- Hex Addr	7ACA	31434
x"00",	-- Hex Addr	7ACB	31435
x"00",	-- Hex Addr	7ACC	31436
x"00",	-- Hex Addr	7ACD	31437
x"00",	-- Hex Addr	7ACE	31438
x"00",	-- Hex Addr	7ACF	31439
x"00",	-- Hex Addr	7AD0	31440
x"00",	-- Hex Addr	7AD1	31441
x"00",	-- Hex Addr	7AD2	31442
x"00",	-- Hex Addr	7AD3	31443
x"00",	-- Hex Addr	7AD4	31444
x"00",	-- Hex Addr	7AD5	31445
x"00",	-- Hex Addr	7AD6	31446
x"00",	-- Hex Addr	7AD7	31447
x"00",	-- Hex Addr	7AD8	31448
x"00",	-- Hex Addr	7AD9	31449
x"00",	-- Hex Addr	7ADA	31450
x"00",	-- Hex Addr	7ADB	31451
x"00",	-- Hex Addr	7ADC	31452
x"00",	-- Hex Addr	7ADD	31453
x"00",	-- Hex Addr	7ADE	31454
x"00",	-- Hex Addr	7ADF	31455
x"00",	-- Hex Addr	7AE0	31456
x"00",	-- Hex Addr	7AE1	31457
x"00",	-- Hex Addr	7AE2	31458
x"00",	-- Hex Addr	7AE3	31459
x"00",	-- Hex Addr	7AE4	31460
x"00",	-- Hex Addr	7AE5	31461
x"00",	-- Hex Addr	7AE6	31462
x"00",	-- Hex Addr	7AE7	31463
x"00",	-- Hex Addr	7AE8	31464
x"00",	-- Hex Addr	7AE9	31465
x"00",	-- Hex Addr	7AEA	31466
x"00",	-- Hex Addr	7AEB	31467
x"00",	-- Hex Addr	7AEC	31468
x"00",	-- Hex Addr	7AED	31469
x"00",	-- Hex Addr	7AEE	31470
x"00",	-- Hex Addr	7AEF	31471
x"00",	-- Hex Addr	7AF0	31472
x"00",	-- Hex Addr	7AF1	31473
x"00",	-- Hex Addr	7AF2	31474
x"00",	-- Hex Addr	7AF3	31475
x"00",	-- Hex Addr	7AF4	31476
x"00",	-- Hex Addr	7AF5	31477
x"00",	-- Hex Addr	7AF6	31478
x"00",	-- Hex Addr	7AF7	31479
x"00",	-- Hex Addr	7AF8	31480
x"00",	-- Hex Addr	7AF9	31481
x"00",	-- Hex Addr	7AFA	31482
x"00",	-- Hex Addr	7AFB	31483
x"00",	-- Hex Addr	7AFC	31484
x"00",	-- Hex Addr	7AFD	31485
x"00",	-- Hex Addr	7AFE	31486
x"00",	-- Hex Addr	7AFF	31487
x"00",	-- Hex Addr	7B00	31488
x"00",	-- Hex Addr	7B01	31489
x"00",	-- Hex Addr	7B02	31490
x"00",	-- Hex Addr	7B03	31491
x"00",	-- Hex Addr	7B04	31492
x"00",	-- Hex Addr	7B05	31493
x"00",	-- Hex Addr	7B06	31494
x"00",	-- Hex Addr	7B07	31495
x"00",	-- Hex Addr	7B08	31496
x"00",	-- Hex Addr	7B09	31497
x"00",	-- Hex Addr	7B0A	31498
x"00",	-- Hex Addr	7B0B	31499
x"00",	-- Hex Addr	7B0C	31500
x"00",	-- Hex Addr	7B0D	31501
x"00",	-- Hex Addr	7B0E	31502
x"00",	-- Hex Addr	7B0F	31503
x"00",	-- Hex Addr	7B10	31504
x"00",	-- Hex Addr	7B11	31505
x"00",	-- Hex Addr	7B12	31506
x"00",	-- Hex Addr	7B13	31507
x"00",	-- Hex Addr	7B14	31508
x"00",	-- Hex Addr	7B15	31509
x"00",	-- Hex Addr	7B16	31510
x"00",	-- Hex Addr	7B17	31511
x"00",	-- Hex Addr	7B18	31512
x"00",	-- Hex Addr	7B19	31513
x"00",	-- Hex Addr	7B1A	31514
x"00",	-- Hex Addr	7B1B	31515
x"00",	-- Hex Addr	7B1C	31516
x"00",	-- Hex Addr	7B1D	31517
x"00",	-- Hex Addr	7B1E	31518
x"00",	-- Hex Addr	7B1F	31519
x"00",	-- Hex Addr	7B20	31520
x"00",	-- Hex Addr	7B21	31521
x"00",	-- Hex Addr	7B22	31522
x"00",	-- Hex Addr	7B23	31523
x"00",	-- Hex Addr	7B24	31524
x"00",	-- Hex Addr	7B25	31525
x"00",	-- Hex Addr	7B26	31526
x"00",	-- Hex Addr	7B27	31527
x"00",	-- Hex Addr	7B28	31528
x"00",	-- Hex Addr	7B29	31529
x"00",	-- Hex Addr	7B2A	31530
x"00",	-- Hex Addr	7B2B	31531
x"00",	-- Hex Addr	7B2C	31532
x"00",	-- Hex Addr	7B2D	31533
x"00",	-- Hex Addr	7B2E	31534
x"00",	-- Hex Addr	7B2F	31535
x"00",	-- Hex Addr	7B30	31536
x"00",	-- Hex Addr	7B31	31537
x"00",	-- Hex Addr	7B32	31538
x"00",	-- Hex Addr	7B33	31539
x"00",	-- Hex Addr	7B34	31540
x"00",	-- Hex Addr	7B35	31541
x"00",	-- Hex Addr	7B36	31542
x"00",	-- Hex Addr	7B37	31543
x"00",	-- Hex Addr	7B38	31544
x"00",	-- Hex Addr	7B39	31545
x"00",	-- Hex Addr	7B3A	31546
x"00",	-- Hex Addr	7B3B	31547
x"00",	-- Hex Addr	7B3C	31548
x"00",	-- Hex Addr	7B3D	31549
x"00",	-- Hex Addr	7B3E	31550
x"00",	-- Hex Addr	7B3F	31551
x"00",	-- Hex Addr	7B40	31552
x"00",	-- Hex Addr	7B41	31553
x"00",	-- Hex Addr	7B42	31554
x"00",	-- Hex Addr	7B43	31555
x"00",	-- Hex Addr	7B44	31556
x"00",	-- Hex Addr	7B45	31557
x"00",	-- Hex Addr	7B46	31558
x"00",	-- Hex Addr	7B47	31559
x"00",	-- Hex Addr	7B48	31560
x"00",	-- Hex Addr	7B49	31561
x"00",	-- Hex Addr	7B4A	31562
x"00",	-- Hex Addr	7B4B	31563
x"00",	-- Hex Addr	7B4C	31564
x"00",	-- Hex Addr	7B4D	31565
x"00",	-- Hex Addr	7B4E	31566
x"00",	-- Hex Addr	7B4F	31567
x"00",	-- Hex Addr	7B50	31568
x"00",	-- Hex Addr	7B51	31569
x"00",	-- Hex Addr	7B52	31570
x"00",	-- Hex Addr	7B53	31571
x"00",	-- Hex Addr	7B54	31572
x"00",	-- Hex Addr	7B55	31573
x"00",	-- Hex Addr	7B56	31574
x"00",	-- Hex Addr	7B57	31575
x"00",	-- Hex Addr	7B58	31576
x"00",	-- Hex Addr	7B59	31577
x"00",	-- Hex Addr	7B5A	31578
x"00",	-- Hex Addr	7B5B	31579
x"00",	-- Hex Addr	7B5C	31580
x"00",	-- Hex Addr	7B5D	31581
x"00",	-- Hex Addr	7B5E	31582
x"00",	-- Hex Addr	7B5F	31583
x"00",	-- Hex Addr	7B60	31584
x"00",	-- Hex Addr	7B61	31585
x"00",	-- Hex Addr	7B62	31586
x"00",	-- Hex Addr	7B63	31587
x"00",	-- Hex Addr	7B64	31588
x"00",	-- Hex Addr	7B65	31589
x"00",	-- Hex Addr	7B66	31590
x"00",	-- Hex Addr	7B67	31591
x"00",	-- Hex Addr	7B68	31592
x"00",	-- Hex Addr	7B69	31593
x"00",	-- Hex Addr	7B6A	31594
x"00",	-- Hex Addr	7B6B	31595
x"00",	-- Hex Addr	7B6C	31596
x"00",	-- Hex Addr	7B6D	31597
x"00",	-- Hex Addr	7B6E	31598
x"00",	-- Hex Addr	7B6F	31599
x"00",	-- Hex Addr	7B70	31600
x"00",	-- Hex Addr	7B71	31601
x"00",	-- Hex Addr	7B72	31602
x"00",	-- Hex Addr	7B73	31603
x"00",	-- Hex Addr	7B74	31604
x"00",	-- Hex Addr	7B75	31605
x"00",	-- Hex Addr	7B76	31606
x"00",	-- Hex Addr	7B77	31607
x"00",	-- Hex Addr	7B78	31608
x"00",	-- Hex Addr	7B79	31609
x"00",	-- Hex Addr	7B7A	31610
x"00",	-- Hex Addr	7B7B	31611
x"00",	-- Hex Addr	7B7C	31612
x"00",	-- Hex Addr	7B7D	31613
x"00",	-- Hex Addr	7B7E	31614
x"00",	-- Hex Addr	7B7F	31615
x"00",	-- Hex Addr	7B80	31616
x"00",	-- Hex Addr	7B81	31617
x"00",	-- Hex Addr	7B82	31618
x"00",	-- Hex Addr	7B83	31619
x"00",	-- Hex Addr	7B84	31620
x"00",	-- Hex Addr	7B85	31621
x"00",	-- Hex Addr	7B86	31622
x"00",	-- Hex Addr	7B87	31623
x"00",	-- Hex Addr	7B88	31624
x"00",	-- Hex Addr	7B89	31625
x"00",	-- Hex Addr	7B8A	31626
x"00",	-- Hex Addr	7B8B	31627
x"00",	-- Hex Addr	7B8C	31628
x"00",	-- Hex Addr	7B8D	31629
x"00",	-- Hex Addr	7B8E	31630
x"00",	-- Hex Addr	7B8F	31631
x"00",	-- Hex Addr	7B90	31632
x"00",	-- Hex Addr	7B91	31633
x"00",	-- Hex Addr	7B92	31634
x"00",	-- Hex Addr	7B93	31635
x"00",	-- Hex Addr	7B94	31636
x"00",	-- Hex Addr	7B95	31637
x"00",	-- Hex Addr	7B96	31638
x"00",	-- Hex Addr	7B97	31639
x"00",	-- Hex Addr	7B98	31640
x"00",	-- Hex Addr	7B99	31641
x"00",	-- Hex Addr	7B9A	31642
x"00",	-- Hex Addr	7B9B	31643
x"00",	-- Hex Addr	7B9C	31644
x"00",	-- Hex Addr	7B9D	31645
x"00",	-- Hex Addr	7B9E	31646
x"00",	-- Hex Addr	7B9F	31647
x"00",	-- Hex Addr	7BA0	31648
x"00",	-- Hex Addr	7BA1	31649
x"00",	-- Hex Addr	7BA2	31650
x"00",	-- Hex Addr	7BA3	31651
x"00",	-- Hex Addr	7BA4	31652
x"00",	-- Hex Addr	7BA5	31653
x"00",	-- Hex Addr	7BA6	31654
x"00",	-- Hex Addr	7BA7	31655
x"00",	-- Hex Addr	7BA8	31656
x"00",	-- Hex Addr	7BA9	31657
x"00",	-- Hex Addr	7BAA	31658
x"00",	-- Hex Addr	7BAB	31659
x"00",	-- Hex Addr	7BAC	31660
x"00",	-- Hex Addr	7BAD	31661
x"00",	-- Hex Addr	7BAE	31662
x"00",	-- Hex Addr	7BAF	31663
x"00",	-- Hex Addr	7BB0	31664
x"00",	-- Hex Addr	7BB1	31665
x"00",	-- Hex Addr	7BB2	31666
x"00",	-- Hex Addr	7BB3	31667
x"00",	-- Hex Addr	7BB4	31668
x"00",	-- Hex Addr	7BB5	31669
x"00",	-- Hex Addr	7BB6	31670
x"00",	-- Hex Addr	7BB7	31671
x"00",	-- Hex Addr	7BB8	31672
x"00",	-- Hex Addr	7BB9	31673
x"00",	-- Hex Addr	7BBA	31674
x"00",	-- Hex Addr	7BBB	31675
x"00",	-- Hex Addr	7BBC	31676
x"00",	-- Hex Addr	7BBD	31677
x"00",	-- Hex Addr	7BBE	31678
x"00",	-- Hex Addr	7BBF	31679
x"00",	-- Hex Addr	7BC0	31680
x"00",	-- Hex Addr	7BC1	31681
x"00",	-- Hex Addr	7BC2	31682
x"00",	-- Hex Addr	7BC3	31683
x"00",	-- Hex Addr	7BC4	31684
x"00",	-- Hex Addr	7BC5	31685
x"00",	-- Hex Addr	7BC6	31686
x"00",	-- Hex Addr	7BC7	31687
x"00",	-- Hex Addr	7BC8	31688
x"00",	-- Hex Addr	7BC9	31689
x"00",	-- Hex Addr	7BCA	31690
x"00",	-- Hex Addr	7BCB	31691
x"00",	-- Hex Addr	7BCC	31692
x"00",	-- Hex Addr	7BCD	31693
x"00",	-- Hex Addr	7BCE	31694
x"00",	-- Hex Addr	7BCF	31695
x"00",	-- Hex Addr	7BD0	31696
x"00",	-- Hex Addr	7BD1	31697
x"00",	-- Hex Addr	7BD2	31698
x"00",	-- Hex Addr	7BD3	31699
x"00",	-- Hex Addr	7BD4	31700
x"00",	-- Hex Addr	7BD5	31701
x"00",	-- Hex Addr	7BD6	31702
x"00",	-- Hex Addr	7BD7	31703
x"00",	-- Hex Addr	7BD8	31704
x"00",	-- Hex Addr	7BD9	31705
x"00",	-- Hex Addr	7BDA	31706
x"00",	-- Hex Addr	7BDB	31707
x"00",	-- Hex Addr	7BDC	31708
x"00",	-- Hex Addr	7BDD	31709
x"00",	-- Hex Addr	7BDE	31710
x"00",	-- Hex Addr	7BDF	31711
x"00",	-- Hex Addr	7BE0	31712
x"00",	-- Hex Addr	7BE1	31713
x"00",	-- Hex Addr	7BE2	31714
x"00",	-- Hex Addr	7BE3	31715
x"00",	-- Hex Addr	7BE4	31716
x"00",	-- Hex Addr	7BE5	31717
x"00",	-- Hex Addr	7BE6	31718
x"00",	-- Hex Addr	7BE7	31719
x"00",	-- Hex Addr	7BE8	31720
x"00",	-- Hex Addr	7BE9	31721
x"00",	-- Hex Addr	7BEA	31722
x"00",	-- Hex Addr	7BEB	31723
x"00",	-- Hex Addr	7BEC	31724
x"00",	-- Hex Addr	7BED	31725
x"00",	-- Hex Addr	7BEE	31726
x"00",	-- Hex Addr	7BEF	31727
x"00",	-- Hex Addr	7BF0	31728
x"00",	-- Hex Addr	7BF1	31729
x"00",	-- Hex Addr	7BF2	31730
x"00",	-- Hex Addr	7BF3	31731
x"00",	-- Hex Addr	7BF4	31732
x"00",	-- Hex Addr	7BF5	31733
x"00",	-- Hex Addr	7BF6	31734
x"00",	-- Hex Addr	7BF7	31735
x"00",	-- Hex Addr	7BF8	31736
x"00",	-- Hex Addr	7BF9	31737
x"00",	-- Hex Addr	7BFA	31738
x"00",	-- Hex Addr	7BFB	31739
x"00",	-- Hex Addr	7BFC	31740
x"00",	-- Hex Addr	7BFD	31741
x"00",	-- Hex Addr	7BFE	31742
x"00",	-- Hex Addr	7BFF	31743
x"00",	-- Hex Addr	7C00	31744
x"00",	-- Hex Addr	7C01	31745
x"00",	-- Hex Addr	7C02	31746
x"00",	-- Hex Addr	7C03	31747
x"00",	-- Hex Addr	7C04	31748
x"00",	-- Hex Addr	7C05	31749
x"00",	-- Hex Addr	7C06	31750
x"00",	-- Hex Addr	7C07	31751
x"00",	-- Hex Addr	7C08	31752
x"00",	-- Hex Addr	7C09	31753
x"00",	-- Hex Addr	7C0A	31754
x"00",	-- Hex Addr	7C0B	31755
x"00",	-- Hex Addr	7C0C	31756
x"00",	-- Hex Addr	7C0D	31757
x"00",	-- Hex Addr	7C0E	31758
x"00",	-- Hex Addr	7C0F	31759
x"00",	-- Hex Addr	7C10	31760
x"00",	-- Hex Addr	7C11	31761
x"00",	-- Hex Addr	7C12	31762
x"00",	-- Hex Addr	7C13	31763
x"00",	-- Hex Addr	7C14	31764
x"00",	-- Hex Addr	7C15	31765
x"00",	-- Hex Addr	7C16	31766
x"00",	-- Hex Addr	7C17	31767
x"00",	-- Hex Addr	7C18	31768
x"00",	-- Hex Addr	7C19	31769
x"00",	-- Hex Addr	7C1A	31770
x"00",	-- Hex Addr	7C1B	31771
x"00",	-- Hex Addr	7C1C	31772
x"00",	-- Hex Addr	7C1D	31773
x"00",	-- Hex Addr	7C1E	31774
x"00",	-- Hex Addr	7C1F	31775
x"00",	-- Hex Addr	7C20	31776
x"00",	-- Hex Addr	7C21	31777
x"00",	-- Hex Addr	7C22	31778
x"00",	-- Hex Addr	7C23	31779
x"00",	-- Hex Addr	7C24	31780
x"00",	-- Hex Addr	7C25	31781
x"00",	-- Hex Addr	7C26	31782
x"00",	-- Hex Addr	7C27	31783
x"00",	-- Hex Addr	7C28	31784
x"00",	-- Hex Addr	7C29	31785
x"00",	-- Hex Addr	7C2A	31786
x"00",	-- Hex Addr	7C2B	31787
x"00",	-- Hex Addr	7C2C	31788
x"00",	-- Hex Addr	7C2D	31789
x"00",	-- Hex Addr	7C2E	31790
x"00",	-- Hex Addr	7C2F	31791
x"00",	-- Hex Addr	7C30	31792
x"00",	-- Hex Addr	7C31	31793
x"00",	-- Hex Addr	7C32	31794
x"00",	-- Hex Addr	7C33	31795
x"00",	-- Hex Addr	7C34	31796
x"00",	-- Hex Addr	7C35	31797
x"00",	-- Hex Addr	7C36	31798
x"00",	-- Hex Addr	7C37	31799
x"00",	-- Hex Addr	7C38	31800
x"00",	-- Hex Addr	7C39	31801
x"00",	-- Hex Addr	7C3A	31802
x"00",	-- Hex Addr	7C3B	31803
x"00",	-- Hex Addr	7C3C	31804
x"00",	-- Hex Addr	7C3D	31805
x"00",	-- Hex Addr	7C3E	31806
x"00",	-- Hex Addr	7C3F	31807
x"00",	-- Hex Addr	7C40	31808
x"00",	-- Hex Addr	7C41	31809
x"00",	-- Hex Addr	7C42	31810
x"00",	-- Hex Addr	7C43	31811
x"00",	-- Hex Addr	7C44	31812
x"00",	-- Hex Addr	7C45	31813
x"00",	-- Hex Addr	7C46	31814
x"00",	-- Hex Addr	7C47	31815
x"00",	-- Hex Addr	7C48	31816
x"00",	-- Hex Addr	7C49	31817
x"00",	-- Hex Addr	7C4A	31818
x"00",	-- Hex Addr	7C4B	31819
x"00",	-- Hex Addr	7C4C	31820
x"00",	-- Hex Addr	7C4D	31821
x"00",	-- Hex Addr	7C4E	31822
x"00",	-- Hex Addr	7C4F	31823
x"00",	-- Hex Addr	7C50	31824
x"00",	-- Hex Addr	7C51	31825
x"00",	-- Hex Addr	7C52	31826
x"00",	-- Hex Addr	7C53	31827
x"00",	-- Hex Addr	7C54	31828
x"00",	-- Hex Addr	7C55	31829
x"00",	-- Hex Addr	7C56	31830
x"00",	-- Hex Addr	7C57	31831
x"00",	-- Hex Addr	7C58	31832
x"00",	-- Hex Addr	7C59	31833
x"00",	-- Hex Addr	7C5A	31834
x"00",	-- Hex Addr	7C5B	31835
x"00",	-- Hex Addr	7C5C	31836
x"00",	-- Hex Addr	7C5D	31837
x"00",	-- Hex Addr	7C5E	31838
x"00",	-- Hex Addr	7C5F	31839
x"00",	-- Hex Addr	7C60	31840
x"00",	-- Hex Addr	7C61	31841
x"00",	-- Hex Addr	7C62	31842
x"00",	-- Hex Addr	7C63	31843
x"00",	-- Hex Addr	7C64	31844
x"00",	-- Hex Addr	7C65	31845
x"00",	-- Hex Addr	7C66	31846
x"00",	-- Hex Addr	7C67	31847
x"00",	-- Hex Addr	7C68	31848
x"00",	-- Hex Addr	7C69	31849
x"00",	-- Hex Addr	7C6A	31850
x"00",	-- Hex Addr	7C6B	31851
x"00",	-- Hex Addr	7C6C	31852
x"00",	-- Hex Addr	7C6D	31853
x"00",	-- Hex Addr	7C6E	31854
x"00",	-- Hex Addr	7C6F	31855
x"00",	-- Hex Addr	7C70	31856
x"00",	-- Hex Addr	7C71	31857
x"00",	-- Hex Addr	7C72	31858
x"00",	-- Hex Addr	7C73	31859
x"00",	-- Hex Addr	7C74	31860
x"00",	-- Hex Addr	7C75	31861
x"00",	-- Hex Addr	7C76	31862
x"00",	-- Hex Addr	7C77	31863
x"00",	-- Hex Addr	7C78	31864
x"00",	-- Hex Addr	7C79	31865
x"00",	-- Hex Addr	7C7A	31866
x"00",	-- Hex Addr	7C7B	31867
x"00",	-- Hex Addr	7C7C	31868
x"00",	-- Hex Addr	7C7D	31869
x"00",	-- Hex Addr	7C7E	31870
x"00",	-- Hex Addr	7C7F	31871
x"00",	-- Hex Addr	7C80	31872
x"00",	-- Hex Addr	7C81	31873
x"00",	-- Hex Addr	7C82	31874
x"00",	-- Hex Addr	7C83	31875
x"00",	-- Hex Addr	7C84	31876
x"00",	-- Hex Addr	7C85	31877
x"00",	-- Hex Addr	7C86	31878
x"00",	-- Hex Addr	7C87	31879
x"00",	-- Hex Addr	7C88	31880
x"00",	-- Hex Addr	7C89	31881
x"00",	-- Hex Addr	7C8A	31882
x"00",	-- Hex Addr	7C8B	31883
x"00",	-- Hex Addr	7C8C	31884
x"00",	-- Hex Addr	7C8D	31885
x"00",	-- Hex Addr	7C8E	31886
x"00",	-- Hex Addr	7C8F	31887
x"00",	-- Hex Addr	7C90	31888
x"00",	-- Hex Addr	7C91	31889
x"00",	-- Hex Addr	7C92	31890
x"00",	-- Hex Addr	7C93	31891
x"00",	-- Hex Addr	7C94	31892
x"00",	-- Hex Addr	7C95	31893
x"00",	-- Hex Addr	7C96	31894
x"00",	-- Hex Addr	7C97	31895
x"00",	-- Hex Addr	7C98	31896
x"00",	-- Hex Addr	7C99	31897
x"00",	-- Hex Addr	7C9A	31898
x"00",	-- Hex Addr	7C9B	31899
x"00",	-- Hex Addr	7C9C	31900
x"00",	-- Hex Addr	7C9D	31901
x"00",	-- Hex Addr	7C9E	31902
x"00",	-- Hex Addr	7C9F	31903
x"00",	-- Hex Addr	7CA0	31904
x"00",	-- Hex Addr	7CA1	31905
x"00",	-- Hex Addr	7CA2	31906
x"00",	-- Hex Addr	7CA3	31907
x"00",	-- Hex Addr	7CA4	31908
x"00",	-- Hex Addr	7CA5	31909
x"00",	-- Hex Addr	7CA6	31910
x"00",	-- Hex Addr	7CA7	31911
x"00",	-- Hex Addr	7CA8	31912
x"00",	-- Hex Addr	7CA9	31913
x"00",	-- Hex Addr	7CAA	31914
x"00",	-- Hex Addr	7CAB	31915
x"00",	-- Hex Addr	7CAC	31916
x"00",	-- Hex Addr	7CAD	31917
x"00",	-- Hex Addr	7CAE	31918
x"00",	-- Hex Addr	7CAF	31919
x"00",	-- Hex Addr	7CB0	31920
x"00",	-- Hex Addr	7CB1	31921
x"00",	-- Hex Addr	7CB2	31922
x"00",	-- Hex Addr	7CB3	31923
x"00",	-- Hex Addr	7CB4	31924
x"00",	-- Hex Addr	7CB5	31925
x"00",	-- Hex Addr	7CB6	31926
x"00",	-- Hex Addr	7CB7	31927
x"00",	-- Hex Addr	7CB8	31928
x"00",	-- Hex Addr	7CB9	31929
x"00",	-- Hex Addr	7CBA	31930
x"00",	-- Hex Addr	7CBB	31931
x"00",	-- Hex Addr	7CBC	31932
x"00",	-- Hex Addr	7CBD	31933
x"00",	-- Hex Addr	7CBE	31934
x"00",	-- Hex Addr	7CBF	31935
x"00",	-- Hex Addr	7CC0	31936
x"00",	-- Hex Addr	7CC1	31937
x"00",	-- Hex Addr	7CC2	31938
x"00",	-- Hex Addr	7CC3	31939
x"00",	-- Hex Addr	7CC4	31940
x"00",	-- Hex Addr	7CC5	31941
x"00",	-- Hex Addr	7CC6	31942
x"00",	-- Hex Addr	7CC7	31943
x"00",	-- Hex Addr	7CC8	31944
x"00",	-- Hex Addr	7CC9	31945
x"00",	-- Hex Addr	7CCA	31946
x"00",	-- Hex Addr	7CCB	31947
x"00",	-- Hex Addr	7CCC	31948
x"00",	-- Hex Addr	7CCD	31949
x"00",	-- Hex Addr	7CCE	31950
x"00",	-- Hex Addr	7CCF	31951
x"00",	-- Hex Addr	7CD0	31952
x"00",	-- Hex Addr	7CD1	31953
x"00",	-- Hex Addr	7CD2	31954
x"00",	-- Hex Addr	7CD3	31955
x"00",	-- Hex Addr	7CD4	31956
x"00",	-- Hex Addr	7CD5	31957
x"00",	-- Hex Addr	7CD6	31958
x"00",	-- Hex Addr	7CD7	31959
x"00",	-- Hex Addr	7CD8	31960
x"00",	-- Hex Addr	7CD9	31961
x"00",	-- Hex Addr	7CDA	31962
x"00",	-- Hex Addr	7CDB	31963
x"00",	-- Hex Addr	7CDC	31964
x"00",	-- Hex Addr	7CDD	31965
x"00",	-- Hex Addr	7CDE	31966
x"00",	-- Hex Addr	7CDF	31967
x"00",	-- Hex Addr	7CE0	31968
x"00",	-- Hex Addr	7CE1	31969
x"00",	-- Hex Addr	7CE2	31970
x"00",	-- Hex Addr	7CE3	31971
x"00",	-- Hex Addr	7CE4	31972
x"00",	-- Hex Addr	7CE5	31973
x"00",	-- Hex Addr	7CE6	31974
x"00",	-- Hex Addr	7CE7	31975
x"00",	-- Hex Addr	7CE8	31976
x"00",	-- Hex Addr	7CE9	31977
x"00",	-- Hex Addr	7CEA	31978
x"00",	-- Hex Addr	7CEB	31979
x"00",	-- Hex Addr	7CEC	31980
x"00",	-- Hex Addr	7CED	31981
x"00",	-- Hex Addr	7CEE	31982
x"00",	-- Hex Addr	7CEF	31983
x"00",	-- Hex Addr	7CF0	31984
x"00",	-- Hex Addr	7CF1	31985
x"00",	-- Hex Addr	7CF2	31986
x"00",	-- Hex Addr	7CF3	31987
x"00",	-- Hex Addr	7CF4	31988
x"00",	-- Hex Addr	7CF5	31989
x"00",	-- Hex Addr	7CF6	31990
x"00",	-- Hex Addr	7CF7	31991
x"00",	-- Hex Addr	7CF8	31992
x"00",	-- Hex Addr	7CF9	31993
x"00",	-- Hex Addr	7CFA	31994
x"00",	-- Hex Addr	7CFB	31995
x"00",	-- Hex Addr	7CFC	31996
x"00",	-- Hex Addr	7CFD	31997
x"00",	-- Hex Addr	7CFE	31998
x"00",	-- Hex Addr	7CFF	31999
x"00",	-- Hex Addr	7D00	32000
x"00",	-- Hex Addr	7D01	32001
x"00",	-- Hex Addr	7D02	32002
x"00",	-- Hex Addr	7D03	32003
x"00",	-- Hex Addr	7D04	32004
x"00",	-- Hex Addr	7D05	32005
x"00",	-- Hex Addr	7D06	32006
x"00",	-- Hex Addr	7D07	32007
x"00",	-- Hex Addr	7D08	32008
x"00",	-- Hex Addr	7D09	32009
x"00",	-- Hex Addr	7D0A	32010
x"00",	-- Hex Addr	7D0B	32011
x"00",	-- Hex Addr	7D0C	32012
x"00",	-- Hex Addr	7D0D	32013
x"00",	-- Hex Addr	7D0E	32014
x"00",	-- Hex Addr	7D0F	32015
x"00",	-- Hex Addr	7D10	32016
x"00",	-- Hex Addr	7D11	32017
x"00",	-- Hex Addr	7D12	32018
x"00",	-- Hex Addr	7D13	32019
x"00",	-- Hex Addr	7D14	32020
x"00",	-- Hex Addr	7D15	32021
x"00",	-- Hex Addr	7D16	32022
x"00",	-- Hex Addr	7D17	32023
x"00",	-- Hex Addr	7D18	32024
x"00",	-- Hex Addr	7D19	32025
x"00",	-- Hex Addr	7D1A	32026
x"00",	-- Hex Addr	7D1B	32027
x"00",	-- Hex Addr	7D1C	32028
x"00",	-- Hex Addr	7D1D	32029
x"00",	-- Hex Addr	7D1E	32030
x"00",	-- Hex Addr	7D1F	32031
x"00",	-- Hex Addr	7D20	32032
x"00",	-- Hex Addr	7D21	32033
x"00",	-- Hex Addr	7D22	32034
x"00",	-- Hex Addr	7D23	32035
x"00",	-- Hex Addr	7D24	32036
x"00",	-- Hex Addr	7D25	32037
x"00",	-- Hex Addr	7D26	32038
x"00",	-- Hex Addr	7D27	32039
x"00",	-- Hex Addr	7D28	32040
x"00",	-- Hex Addr	7D29	32041
x"00",	-- Hex Addr	7D2A	32042
x"00",	-- Hex Addr	7D2B	32043
x"00",	-- Hex Addr	7D2C	32044
x"00",	-- Hex Addr	7D2D	32045
x"00",	-- Hex Addr	7D2E	32046
x"00",	-- Hex Addr	7D2F	32047
x"00",	-- Hex Addr	7D30	32048
x"00",	-- Hex Addr	7D31	32049
x"00",	-- Hex Addr	7D32	32050
x"00",	-- Hex Addr	7D33	32051
x"00",	-- Hex Addr	7D34	32052
x"00",	-- Hex Addr	7D35	32053
x"00",	-- Hex Addr	7D36	32054
x"00",	-- Hex Addr	7D37	32055
x"00",	-- Hex Addr	7D38	32056
x"00",	-- Hex Addr	7D39	32057
x"00",	-- Hex Addr	7D3A	32058
x"00",	-- Hex Addr	7D3B	32059
x"00",	-- Hex Addr	7D3C	32060
x"00",	-- Hex Addr	7D3D	32061
x"00",	-- Hex Addr	7D3E	32062
x"00",	-- Hex Addr	7D3F	32063
x"00",	-- Hex Addr	7D40	32064
x"00",	-- Hex Addr	7D41	32065
x"00",	-- Hex Addr	7D42	32066
x"00",	-- Hex Addr	7D43	32067
x"00",	-- Hex Addr	7D44	32068
x"00",	-- Hex Addr	7D45	32069
x"00",	-- Hex Addr	7D46	32070
x"00",	-- Hex Addr	7D47	32071
x"00",	-- Hex Addr	7D48	32072
x"00",	-- Hex Addr	7D49	32073
x"00",	-- Hex Addr	7D4A	32074
x"00",	-- Hex Addr	7D4B	32075
x"00",	-- Hex Addr	7D4C	32076
x"00",	-- Hex Addr	7D4D	32077
x"00",	-- Hex Addr	7D4E	32078
x"00",	-- Hex Addr	7D4F	32079
x"00",	-- Hex Addr	7D50	32080
x"00",	-- Hex Addr	7D51	32081
x"00",	-- Hex Addr	7D52	32082
x"00",	-- Hex Addr	7D53	32083
x"00",	-- Hex Addr	7D54	32084
x"00",	-- Hex Addr	7D55	32085
x"00",	-- Hex Addr	7D56	32086
x"00",	-- Hex Addr	7D57	32087
x"00",	-- Hex Addr	7D58	32088
x"00",	-- Hex Addr	7D59	32089
x"00",	-- Hex Addr	7D5A	32090
x"00",	-- Hex Addr	7D5B	32091
x"00",	-- Hex Addr	7D5C	32092
x"00",	-- Hex Addr	7D5D	32093
x"00",	-- Hex Addr	7D5E	32094
x"00",	-- Hex Addr	7D5F	32095
x"00",	-- Hex Addr	7D60	32096
x"00",	-- Hex Addr	7D61	32097
x"00",	-- Hex Addr	7D62	32098
x"00",	-- Hex Addr	7D63	32099
x"00",	-- Hex Addr	7D64	32100
x"00",	-- Hex Addr	7D65	32101
x"00",	-- Hex Addr	7D66	32102
x"00",	-- Hex Addr	7D67	32103
x"00",	-- Hex Addr	7D68	32104
x"00",	-- Hex Addr	7D69	32105
x"00",	-- Hex Addr	7D6A	32106
x"00",	-- Hex Addr	7D6B	32107
x"00",	-- Hex Addr	7D6C	32108
x"00",	-- Hex Addr	7D6D	32109
x"00",	-- Hex Addr	7D6E	32110
x"00",	-- Hex Addr	7D6F	32111
x"00",	-- Hex Addr	7D70	32112
x"00",	-- Hex Addr	7D71	32113
x"00",	-- Hex Addr	7D72	32114
x"00",	-- Hex Addr	7D73	32115
x"00",	-- Hex Addr	7D74	32116
x"00",	-- Hex Addr	7D75	32117
x"00",	-- Hex Addr	7D76	32118
x"00",	-- Hex Addr	7D77	32119
x"00",	-- Hex Addr	7D78	32120
x"00",	-- Hex Addr	7D79	32121
x"00",	-- Hex Addr	7D7A	32122
x"00",	-- Hex Addr	7D7B	32123
x"00",	-- Hex Addr	7D7C	32124
x"00",	-- Hex Addr	7D7D	32125
x"00",	-- Hex Addr	7D7E	32126
x"00",	-- Hex Addr	7D7F	32127
x"00",	-- Hex Addr	7D80	32128
x"00",	-- Hex Addr	7D81	32129
x"00",	-- Hex Addr	7D82	32130
x"00",	-- Hex Addr	7D83	32131
x"00",	-- Hex Addr	7D84	32132
x"00",	-- Hex Addr	7D85	32133
x"00",	-- Hex Addr	7D86	32134
x"00",	-- Hex Addr	7D87	32135
x"00",	-- Hex Addr	7D88	32136
x"00",	-- Hex Addr	7D89	32137
x"00",	-- Hex Addr	7D8A	32138
x"00",	-- Hex Addr	7D8B	32139
x"00",	-- Hex Addr	7D8C	32140
x"00",	-- Hex Addr	7D8D	32141
x"00",	-- Hex Addr	7D8E	32142
x"00",	-- Hex Addr	7D8F	32143
x"00",	-- Hex Addr	7D90	32144
x"00",	-- Hex Addr	7D91	32145
x"00",	-- Hex Addr	7D92	32146
x"00",	-- Hex Addr	7D93	32147
x"00",	-- Hex Addr	7D94	32148
x"00",	-- Hex Addr	7D95	32149
x"00",	-- Hex Addr	7D96	32150
x"00",	-- Hex Addr	7D97	32151
x"00",	-- Hex Addr	7D98	32152
x"00",	-- Hex Addr	7D99	32153
x"00",	-- Hex Addr	7D9A	32154
x"00",	-- Hex Addr	7D9B	32155
x"00",	-- Hex Addr	7D9C	32156
x"00",	-- Hex Addr	7D9D	32157
x"00",	-- Hex Addr	7D9E	32158
x"00",	-- Hex Addr	7D9F	32159
x"00",	-- Hex Addr	7DA0	32160
x"00",	-- Hex Addr	7DA1	32161
x"00",	-- Hex Addr	7DA2	32162
x"00",	-- Hex Addr	7DA3	32163
x"00",	-- Hex Addr	7DA4	32164
x"00",	-- Hex Addr	7DA5	32165
x"00",	-- Hex Addr	7DA6	32166
x"00",	-- Hex Addr	7DA7	32167
x"00",	-- Hex Addr	7DA8	32168
x"00",	-- Hex Addr	7DA9	32169
x"00",	-- Hex Addr	7DAA	32170
x"00",	-- Hex Addr	7DAB	32171
x"00",	-- Hex Addr	7DAC	32172
x"00",	-- Hex Addr	7DAD	32173
x"00",	-- Hex Addr	7DAE	32174
x"00",	-- Hex Addr	7DAF	32175
x"00",	-- Hex Addr	7DB0	32176
x"00",	-- Hex Addr	7DB1	32177
x"00",	-- Hex Addr	7DB2	32178
x"00",	-- Hex Addr	7DB3	32179
x"00",	-- Hex Addr	7DB4	32180
x"00",	-- Hex Addr	7DB5	32181
x"00",	-- Hex Addr	7DB6	32182
x"00",	-- Hex Addr	7DB7	32183
x"00",	-- Hex Addr	7DB8	32184
x"00",	-- Hex Addr	7DB9	32185
x"00",	-- Hex Addr	7DBA	32186
x"00",	-- Hex Addr	7DBB	32187
x"00",	-- Hex Addr	7DBC	32188
x"00",	-- Hex Addr	7DBD	32189
x"00",	-- Hex Addr	7DBE	32190
x"00",	-- Hex Addr	7DBF	32191
x"00",	-- Hex Addr	7DC0	32192
x"00",	-- Hex Addr	7DC1	32193
x"00",	-- Hex Addr	7DC2	32194
x"00",	-- Hex Addr	7DC3	32195
x"00",	-- Hex Addr	7DC4	32196
x"00",	-- Hex Addr	7DC5	32197
x"00",	-- Hex Addr	7DC6	32198
x"00",	-- Hex Addr	7DC7	32199
x"00",	-- Hex Addr	7DC8	32200
x"00",	-- Hex Addr	7DC9	32201
x"00",	-- Hex Addr	7DCA	32202
x"00",	-- Hex Addr	7DCB	32203
x"00",	-- Hex Addr	7DCC	32204
x"00",	-- Hex Addr	7DCD	32205
x"00",	-- Hex Addr	7DCE	32206
x"00",	-- Hex Addr	7DCF	32207
x"00",	-- Hex Addr	7DD0	32208
x"00",	-- Hex Addr	7DD1	32209
x"00",	-- Hex Addr	7DD2	32210
x"00",	-- Hex Addr	7DD3	32211
x"00",	-- Hex Addr	7DD4	32212
x"00",	-- Hex Addr	7DD5	32213
x"00",	-- Hex Addr	7DD6	32214
x"00",	-- Hex Addr	7DD7	32215
x"00",	-- Hex Addr	7DD8	32216
x"00",	-- Hex Addr	7DD9	32217
x"00",	-- Hex Addr	7DDA	32218
x"00",	-- Hex Addr	7DDB	32219
x"00",	-- Hex Addr	7DDC	32220
x"00",	-- Hex Addr	7DDD	32221
x"00",	-- Hex Addr	7DDE	32222
x"00",	-- Hex Addr	7DDF	32223
x"00",	-- Hex Addr	7DE0	32224
x"00",	-- Hex Addr	7DE1	32225
x"00",	-- Hex Addr	7DE2	32226
x"00",	-- Hex Addr	7DE3	32227
x"00",	-- Hex Addr	7DE4	32228
x"00",	-- Hex Addr	7DE5	32229
x"00",	-- Hex Addr	7DE6	32230
x"00",	-- Hex Addr	7DE7	32231
x"00",	-- Hex Addr	7DE8	32232
x"00",	-- Hex Addr	7DE9	32233
x"00",	-- Hex Addr	7DEA	32234
x"00",	-- Hex Addr	7DEB	32235
x"00",	-- Hex Addr	7DEC	32236
x"00",	-- Hex Addr	7DED	32237
x"00",	-- Hex Addr	7DEE	32238
x"00",	-- Hex Addr	7DEF	32239
x"00",	-- Hex Addr	7DF0	32240
x"00",	-- Hex Addr	7DF1	32241
x"00",	-- Hex Addr	7DF2	32242
x"00",	-- Hex Addr	7DF3	32243
x"00",	-- Hex Addr	7DF4	32244
x"00",	-- Hex Addr	7DF5	32245
x"00",	-- Hex Addr	7DF6	32246
x"00",	-- Hex Addr	7DF7	32247
x"00",	-- Hex Addr	7DF8	32248
x"00",	-- Hex Addr	7DF9	32249
x"00",	-- Hex Addr	7DFA	32250
x"00",	-- Hex Addr	7DFB	32251
x"00",	-- Hex Addr	7DFC	32252
x"00",	-- Hex Addr	7DFD	32253
x"00",	-- Hex Addr	7DFE	32254
x"00",	-- Hex Addr	7DFF	32255
x"00",	-- Hex Addr	7E00	32256
x"00",	-- Hex Addr	7E01	32257
x"00",	-- Hex Addr	7E02	32258
x"00",	-- Hex Addr	7E03	32259
x"00",	-- Hex Addr	7E04	32260
x"00",	-- Hex Addr	7E05	32261
x"00",	-- Hex Addr	7E06	32262
x"00",	-- Hex Addr	7E07	32263
x"00",	-- Hex Addr	7E08	32264
x"00",	-- Hex Addr	7E09	32265
x"00",	-- Hex Addr	7E0A	32266
x"00",	-- Hex Addr	7E0B	32267
x"00",	-- Hex Addr	7E0C	32268
x"00",	-- Hex Addr	7E0D	32269
x"00",	-- Hex Addr	7E0E	32270
x"00",	-- Hex Addr	7E0F	32271
x"00",	-- Hex Addr	7E10	32272
x"00",	-- Hex Addr	7E11	32273
x"00",	-- Hex Addr	7E12	32274
x"00",	-- Hex Addr	7E13	32275
x"00",	-- Hex Addr	7E14	32276
x"00",	-- Hex Addr	7E15	32277
x"00",	-- Hex Addr	7E16	32278
x"00",	-- Hex Addr	7E17	32279
x"00",	-- Hex Addr	7E18	32280
x"00",	-- Hex Addr	7E19	32281
x"00",	-- Hex Addr	7E1A	32282
x"00",	-- Hex Addr	7E1B	32283
x"00",	-- Hex Addr	7E1C	32284
x"00",	-- Hex Addr	7E1D	32285
x"00",	-- Hex Addr	7E1E	32286
x"00",	-- Hex Addr	7E1F	32287
x"00",	-- Hex Addr	7E20	32288
x"00",	-- Hex Addr	7E21	32289
x"00",	-- Hex Addr	7E22	32290
x"00",	-- Hex Addr	7E23	32291
x"00",	-- Hex Addr	7E24	32292
x"00",	-- Hex Addr	7E25	32293
x"00",	-- Hex Addr	7E26	32294
x"00",	-- Hex Addr	7E27	32295
x"00",	-- Hex Addr	7E28	32296
x"00",	-- Hex Addr	7E29	32297
x"00",	-- Hex Addr	7E2A	32298
x"00",	-- Hex Addr	7E2B	32299
x"00",	-- Hex Addr	7E2C	32300
x"00",	-- Hex Addr	7E2D	32301
x"00",	-- Hex Addr	7E2E	32302
x"00",	-- Hex Addr	7E2F	32303
x"00",	-- Hex Addr	7E30	32304
x"00",	-- Hex Addr	7E31	32305
x"00",	-- Hex Addr	7E32	32306
x"00",	-- Hex Addr	7E33	32307
x"00",	-- Hex Addr	7E34	32308
x"00",	-- Hex Addr	7E35	32309
x"00",	-- Hex Addr	7E36	32310
x"00",	-- Hex Addr	7E37	32311
x"00",	-- Hex Addr	7E38	32312
x"00",	-- Hex Addr	7E39	32313
x"00",	-- Hex Addr	7E3A	32314
x"00",	-- Hex Addr	7E3B	32315
x"00",	-- Hex Addr	7E3C	32316
x"00",	-- Hex Addr	7E3D	32317
x"00",	-- Hex Addr	7E3E	32318
x"00",	-- Hex Addr	7E3F	32319
x"00",	-- Hex Addr	7E40	32320
x"00",	-- Hex Addr	7E41	32321
x"00",	-- Hex Addr	7E42	32322
x"00",	-- Hex Addr	7E43	32323
x"00",	-- Hex Addr	7E44	32324
x"00",	-- Hex Addr	7E45	32325
x"00",	-- Hex Addr	7E46	32326
x"00",	-- Hex Addr	7E47	32327
x"00",	-- Hex Addr	7E48	32328
x"00",	-- Hex Addr	7E49	32329
x"00",	-- Hex Addr	7E4A	32330
x"00",	-- Hex Addr	7E4B	32331
x"00",	-- Hex Addr	7E4C	32332
x"00",	-- Hex Addr	7E4D	32333
x"00",	-- Hex Addr	7E4E	32334
x"00",	-- Hex Addr	7E4F	32335
x"00",	-- Hex Addr	7E50	32336
x"00",	-- Hex Addr	7E51	32337
x"00",	-- Hex Addr	7E52	32338
x"00",	-- Hex Addr	7E53	32339
x"00",	-- Hex Addr	7E54	32340
x"00",	-- Hex Addr	7E55	32341
x"00",	-- Hex Addr	7E56	32342
x"00",	-- Hex Addr	7E57	32343
x"00",	-- Hex Addr	7E58	32344
x"00",	-- Hex Addr	7E59	32345
x"00",	-- Hex Addr	7E5A	32346
x"00",	-- Hex Addr	7E5B	32347
x"00",	-- Hex Addr	7E5C	32348
x"00",	-- Hex Addr	7E5D	32349
x"00",	-- Hex Addr	7E5E	32350
x"00",	-- Hex Addr	7E5F	32351
x"00",	-- Hex Addr	7E60	32352
x"00",	-- Hex Addr	7E61	32353
x"00",	-- Hex Addr	7E62	32354
x"00",	-- Hex Addr	7E63	32355
x"00",	-- Hex Addr	7E64	32356
x"00",	-- Hex Addr	7E65	32357
x"00",	-- Hex Addr	7E66	32358
x"00",	-- Hex Addr	7E67	32359
x"00",	-- Hex Addr	7E68	32360
x"00",	-- Hex Addr	7E69	32361
x"00",	-- Hex Addr	7E6A	32362
x"00",	-- Hex Addr	7E6B	32363
x"00",	-- Hex Addr	7E6C	32364
x"00",	-- Hex Addr	7E6D	32365
x"00",	-- Hex Addr	7E6E	32366
x"00",	-- Hex Addr	7E6F	32367
x"00",	-- Hex Addr	7E70	32368
x"00",	-- Hex Addr	7E71	32369
x"00",	-- Hex Addr	7E72	32370
x"00",	-- Hex Addr	7E73	32371
x"00",	-- Hex Addr	7E74	32372
x"00",	-- Hex Addr	7E75	32373
x"00",	-- Hex Addr	7E76	32374
x"00",	-- Hex Addr	7E77	32375
x"00",	-- Hex Addr	7E78	32376
x"00",	-- Hex Addr	7E79	32377
x"00",	-- Hex Addr	7E7A	32378
x"00",	-- Hex Addr	7E7B	32379
x"00",	-- Hex Addr	7E7C	32380
x"00",	-- Hex Addr	7E7D	32381
x"00",	-- Hex Addr	7E7E	32382
x"00",	-- Hex Addr	7E7F	32383
x"00",	-- Hex Addr	7E80	32384
x"00",	-- Hex Addr	7E81	32385
x"00",	-- Hex Addr	7E82	32386
x"00",	-- Hex Addr	7E83	32387
x"00",	-- Hex Addr	7E84	32388
x"00",	-- Hex Addr	7E85	32389
x"00",	-- Hex Addr	7E86	32390
x"00",	-- Hex Addr	7E87	32391
x"00",	-- Hex Addr	7E88	32392
x"00",	-- Hex Addr	7E89	32393
x"00",	-- Hex Addr	7E8A	32394
x"00",	-- Hex Addr	7E8B	32395
x"00",	-- Hex Addr	7E8C	32396
x"00",	-- Hex Addr	7E8D	32397
x"00",	-- Hex Addr	7E8E	32398
x"00",	-- Hex Addr	7E8F	32399
x"00",	-- Hex Addr	7E90	32400
x"00",	-- Hex Addr	7E91	32401
x"00",	-- Hex Addr	7E92	32402
x"00",	-- Hex Addr	7E93	32403
x"00",	-- Hex Addr	7E94	32404
x"00",	-- Hex Addr	7E95	32405
x"00",	-- Hex Addr	7E96	32406
x"00",	-- Hex Addr	7E97	32407
x"00",	-- Hex Addr	7E98	32408
x"00",	-- Hex Addr	7E99	32409
x"00",	-- Hex Addr	7E9A	32410
x"00",	-- Hex Addr	7E9B	32411
x"00",	-- Hex Addr	7E9C	32412
x"00",	-- Hex Addr	7E9D	32413
x"00",	-- Hex Addr	7E9E	32414
x"00",	-- Hex Addr	7E9F	32415
x"00",	-- Hex Addr	7EA0	32416
x"00",	-- Hex Addr	7EA1	32417
x"00",	-- Hex Addr	7EA2	32418
x"00",	-- Hex Addr	7EA3	32419
x"00",	-- Hex Addr	7EA4	32420
x"00",	-- Hex Addr	7EA5	32421
x"00",	-- Hex Addr	7EA6	32422
x"00",	-- Hex Addr	7EA7	32423
x"00",	-- Hex Addr	7EA8	32424
x"00",	-- Hex Addr	7EA9	32425
x"00",	-- Hex Addr	7EAA	32426
x"00",	-- Hex Addr	7EAB	32427
x"00",	-- Hex Addr	7EAC	32428
x"00",	-- Hex Addr	7EAD	32429
x"00",	-- Hex Addr	7EAE	32430
x"00",	-- Hex Addr	7EAF	32431
x"00",	-- Hex Addr	7EB0	32432
x"00",	-- Hex Addr	7EB1	32433
x"00",	-- Hex Addr	7EB2	32434
x"00",	-- Hex Addr	7EB3	32435
x"00",	-- Hex Addr	7EB4	32436
x"00",	-- Hex Addr	7EB5	32437
x"00",	-- Hex Addr	7EB6	32438
x"00",	-- Hex Addr	7EB7	32439
x"00",	-- Hex Addr	7EB8	32440
x"00",	-- Hex Addr	7EB9	32441
x"00",	-- Hex Addr	7EBA	32442
x"00",	-- Hex Addr	7EBB	32443
x"00",	-- Hex Addr	7EBC	32444
x"00",	-- Hex Addr	7EBD	32445
x"00",	-- Hex Addr	7EBE	32446
x"00",	-- Hex Addr	7EBF	32447
x"00",	-- Hex Addr	7EC0	32448
x"00",	-- Hex Addr	7EC1	32449
x"00",	-- Hex Addr	7EC2	32450
x"00",	-- Hex Addr	7EC3	32451
x"00",	-- Hex Addr	7EC4	32452
x"00",	-- Hex Addr	7EC5	32453
x"00",	-- Hex Addr	7EC6	32454
x"00",	-- Hex Addr	7EC7	32455
x"00",	-- Hex Addr	7EC8	32456
x"00",	-- Hex Addr	7EC9	32457
x"00",	-- Hex Addr	7ECA	32458
x"00",	-- Hex Addr	7ECB	32459
x"00",	-- Hex Addr	7ECC	32460
x"00",	-- Hex Addr	7ECD	32461
x"00",	-- Hex Addr	7ECE	32462
x"00",	-- Hex Addr	7ECF	32463
x"00",	-- Hex Addr	7ED0	32464
x"00",	-- Hex Addr	7ED1	32465
x"00",	-- Hex Addr	7ED2	32466
x"00",	-- Hex Addr	7ED3	32467
x"00",	-- Hex Addr	7ED4	32468
x"00",	-- Hex Addr	7ED5	32469
x"00",	-- Hex Addr	7ED6	32470
x"00",	-- Hex Addr	7ED7	32471
x"00",	-- Hex Addr	7ED8	32472
x"00",	-- Hex Addr	7ED9	32473
x"00",	-- Hex Addr	7EDA	32474
x"00",	-- Hex Addr	7EDB	32475
x"00",	-- Hex Addr	7EDC	32476
x"00",	-- Hex Addr	7EDD	32477
x"00",	-- Hex Addr	7EDE	32478
x"00",	-- Hex Addr	7EDF	32479
x"00",	-- Hex Addr	7EE0	32480
x"00",	-- Hex Addr	7EE1	32481
x"00",	-- Hex Addr	7EE2	32482
x"00",	-- Hex Addr	7EE3	32483
x"00",	-- Hex Addr	7EE4	32484
x"00",	-- Hex Addr	7EE5	32485
x"00",	-- Hex Addr	7EE6	32486
x"00",	-- Hex Addr	7EE7	32487
x"00",	-- Hex Addr	7EE8	32488
x"00",	-- Hex Addr	7EE9	32489
x"00",	-- Hex Addr	7EEA	32490
x"00",	-- Hex Addr	7EEB	32491
x"00",	-- Hex Addr	7EEC	32492
x"00",	-- Hex Addr	7EED	32493
x"00",	-- Hex Addr	7EEE	32494
x"00",	-- Hex Addr	7EEF	32495
x"00",	-- Hex Addr	7EF0	32496
x"00",	-- Hex Addr	7EF1	32497
x"00",	-- Hex Addr	7EF2	32498
x"00",	-- Hex Addr	7EF3	32499
x"00",	-- Hex Addr	7EF4	32500
x"00",	-- Hex Addr	7EF5	32501
x"00",	-- Hex Addr	7EF6	32502
x"00",	-- Hex Addr	7EF7	32503
x"00",	-- Hex Addr	7EF8	32504
x"00",	-- Hex Addr	7EF9	32505
x"00",	-- Hex Addr	7EFA	32506
x"00",	-- Hex Addr	7EFB	32507
x"00",	-- Hex Addr	7EFC	32508
x"00",	-- Hex Addr	7EFD	32509
x"00",	-- Hex Addr	7EFE	32510
x"00",	-- Hex Addr	7EFF	32511
x"00",	-- Hex Addr	7F00	32512
x"00",	-- Hex Addr	7F01	32513
x"00",	-- Hex Addr	7F02	32514
x"00",	-- Hex Addr	7F03	32515
x"00",	-- Hex Addr	7F04	32516
x"00",	-- Hex Addr	7F05	32517
x"00",	-- Hex Addr	7F06	32518
x"00",	-- Hex Addr	7F07	32519
x"00",	-- Hex Addr	7F08	32520
x"00",	-- Hex Addr	7F09	32521
x"00",	-- Hex Addr	7F0A	32522
x"00",	-- Hex Addr	7F0B	32523
x"00",	-- Hex Addr	7F0C	32524
x"00",	-- Hex Addr	7F0D	32525
x"00",	-- Hex Addr	7F0E	32526
x"00",	-- Hex Addr	7F0F	32527
x"00",	-- Hex Addr	7F10	32528
x"00",	-- Hex Addr	7F11	32529
x"00",	-- Hex Addr	7F12	32530
x"00",	-- Hex Addr	7F13	32531
x"00",	-- Hex Addr	7F14	32532
x"00",	-- Hex Addr	7F15	32533
x"00",	-- Hex Addr	7F16	32534
x"00",	-- Hex Addr	7F17	32535
x"00",	-- Hex Addr	7F18	32536
x"00",	-- Hex Addr	7F19	32537
x"00",	-- Hex Addr	7F1A	32538
x"00",	-- Hex Addr	7F1B	32539
x"00",	-- Hex Addr	7F1C	32540
x"00",	-- Hex Addr	7F1D	32541
x"00",	-- Hex Addr	7F1E	32542
x"00",	-- Hex Addr	7F1F	32543
x"00",	-- Hex Addr	7F20	32544
x"00",	-- Hex Addr	7F21	32545
x"00",	-- Hex Addr	7F22	32546
x"00",	-- Hex Addr	7F23	32547
x"00",	-- Hex Addr	7F24	32548
x"00",	-- Hex Addr	7F25	32549
x"00",	-- Hex Addr	7F26	32550
x"00",	-- Hex Addr	7F27	32551
x"00",	-- Hex Addr	7F28	32552
x"00",	-- Hex Addr	7F29	32553
x"00",	-- Hex Addr	7F2A	32554
x"00",	-- Hex Addr	7F2B	32555
x"00",	-- Hex Addr	7F2C	32556
x"00",	-- Hex Addr	7F2D	32557
x"00",	-- Hex Addr	7F2E	32558
x"00",	-- Hex Addr	7F2F	32559
x"00",	-- Hex Addr	7F30	32560
x"00",	-- Hex Addr	7F31	32561
x"00",	-- Hex Addr	7F32	32562
x"00",	-- Hex Addr	7F33	32563
x"00",	-- Hex Addr	7F34	32564
x"00",	-- Hex Addr	7F35	32565
x"00",	-- Hex Addr	7F36	32566
x"00",	-- Hex Addr	7F37	32567
x"00",	-- Hex Addr	7F38	32568
x"00",	-- Hex Addr	7F39	32569
x"00",	-- Hex Addr	7F3A	32570
x"00",	-- Hex Addr	7F3B	32571
x"00",	-- Hex Addr	7F3C	32572
x"00",	-- Hex Addr	7F3D	32573
x"00",	-- Hex Addr	7F3E	32574
x"00",	-- Hex Addr	7F3F	32575
x"00",	-- Hex Addr	7F40	32576
x"00",	-- Hex Addr	7F41	32577
x"00",	-- Hex Addr	7F42	32578
x"00",	-- Hex Addr	7F43	32579
x"00",	-- Hex Addr	7F44	32580
x"00",	-- Hex Addr	7F45	32581
x"00",	-- Hex Addr	7F46	32582
x"00",	-- Hex Addr	7F47	32583
x"00",	-- Hex Addr	7F48	32584
x"00",	-- Hex Addr	7F49	32585
x"00",	-- Hex Addr	7F4A	32586
x"00",	-- Hex Addr	7F4B	32587
x"00",	-- Hex Addr	7F4C	32588
x"00",	-- Hex Addr	7F4D	32589
x"00",	-- Hex Addr	7F4E	32590
x"00",	-- Hex Addr	7F4F	32591
x"00",	-- Hex Addr	7F50	32592
x"00",	-- Hex Addr	7F51	32593
x"00",	-- Hex Addr	7F52	32594
x"00",	-- Hex Addr	7F53	32595
x"00",	-- Hex Addr	7F54	32596
x"00",	-- Hex Addr	7F55	32597
x"00",	-- Hex Addr	7F56	32598
x"00",	-- Hex Addr	7F57	32599
x"00",	-- Hex Addr	7F58	32600
x"00",	-- Hex Addr	7F59	32601
x"00",	-- Hex Addr	7F5A	32602
x"00",	-- Hex Addr	7F5B	32603
x"00",	-- Hex Addr	7F5C	32604
x"00",	-- Hex Addr	7F5D	32605
x"00",	-- Hex Addr	7F5E	32606
x"00",	-- Hex Addr	7F5F	32607
x"00",	-- Hex Addr	7F60	32608
x"00",	-- Hex Addr	7F61	32609
x"00",	-- Hex Addr	7F62	32610
x"00",	-- Hex Addr	7F63	32611
x"00",	-- Hex Addr	7F64	32612
x"00",	-- Hex Addr	7F65	32613
x"00",	-- Hex Addr	7F66	32614
x"00",	-- Hex Addr	7F67	32615
x"00",	-- Hex Addr	7F68	32616
x"00",	-- Hex Addr	7F69	32617
x"00",	-- Hex Addr	7F6A	32618
x"00",	-- Hex Addr	7F6B	32619
x"00",	-- Hex Addr	7F6C	32620
x"00",	-- Hex Addr	7F6D	32621
x"00",	-- Hex Addr	7F6E	32622
x"00",	-- Hex Addr	7F6F	32623
x"00",	-- Hex Addr	7F70	32624
x"00",	-- Hex Addr	7F71	32625
x"00",	-- Hex Addr	7F72	32626
x"00",	-- Hex Addr	7F73	32627
x"00",	-- Hex Addr	7F74	32628
x"00",	-- Hex Addr	7F75	32629
x"00",	-- Hex Addr	7F76	32630
x"00",	-- Hex Addr	7F77	32631
x"00",	-- Hex Addr	7F78	32632
x"00",	-- Hex Addr	7F79	32633
x"00",	-- Hex Addr	7F7A	32634
x"00",	-- Hex Addr	7F7B	32635
x"00",	-- Hex Addr	7F7C	32636
x"00",	-- Hex Addr	7F7D	32637
x"00",	-- Hex Addr	7F7E	32638
x"00",	-- Hex Addr	7F7F	32639
x"00",	-- Hex Addr	7F80	32640
x"00",	-- Hex Addr	7F81	32641
x"00",	-- Hex Addr	7F82	32642
x"00",	-- Hex Addr	7F83	32643
x"00",	-- Hex Addr	7F84	32644
x"00",	-- Hex Addr	7F85	32645
x"00",	-- Hex Addr	7F86	32646
x"00",	-- Hex Addr	7F87	32647
x"00",	-- Hex Addr	7F88	32648
x"00",	-- Hex Addr	7F89	32649
x"00",	-- Hex Addr	7F8A	32650
x"00",	-- Hex Addr	7F8B	32651
x"00",	-- Hex Addr	7F8C	32652
x"00",	-- Hex Addr	7F8D	32653
x"00",	-- Hex Addr	7F8E	32654
x"00",	-- Hex Addr	7F8F	32655
x"00",	-- Hex Addr	7F90	32656
x"00",	-- Hex Addr	7F91	32657
x"00",	-- Hex Addr	7F92	32658
x"00",	-- Hex Addr	7F93	32659
x"00",	-- Hex Addr	7F94	32660
x"00",	-- Hex Addr	7F95	32661
x"00",	-- Hex Addr	7F96	32662
x"00",	-- Hex Addr	7F97	32663
x"00",	-- Hex Addr	7F98	32664
x"00",	-- Hex Addr	7F99	32665
x"00",	-- Hex Addr	7F9A	32666
x"00",	-- Hex Addr	7F9B	32667
x"00",	-- Hex Addr	7F9C	32668
x"00",	-- Hex Addr	7F9D	32669
x"00",	-- Hex Addr	7F9E	32670
x"00",	-- Hex Addr	7F9F	32671
x"00",	-- Hex Addr	7FA0	32672
x"00",	-- Hex Addr	7FA1	32673
x"00",	-- Hex Addr	7FA2	32674
x"00",	-- Hex Addr	7FA3	32675
x"00",	-- Hex Addr	7FA4	32676
x"00",	-- Hex Addr	7FA5	32677
x"00",	-- Hex Addr	7FA6	32678
x"00",	-- Hex Addr	7FA7	32679
x"00",	-- Hex Addr	7FA8	32680
x"00",	-- Hex Addr	7FA9	32681
x"00",	-- Hex Addr	7FAA	32682
x"00",	-- Hex Addr	7FAB	32683
x"00",	-- Hex Addr	7FAC	32684
x"00",	-- Hex Addr	7FAD	32685
x"00",	-- Hex Addr	7FAE	32686
x"00",	-- Hex Addr	7FAF	32687
x"00",	-- Hex Addr	7FB0	32688
x"00",	-- Hex Addr	7FB1	32689
x"00",	-- Hex Addr	7FB2	32690
x"00",	-- Hex Addr	7FB3	32691
x"00",	-- Hex Addr	7FB4	32692
x"00",	-- Hex Addr	7FB5	32693
x"00",	-- Hex Addr	7FB6	32694
x"00",	-- Hex Addr	7FB7	32695
x"00",	-- Hex Addr	7FB8	32696
x"00",	-- Hex Addr	7FB9	32697
x"00",	-- Hex Addr	7FBA	32698
x"00",	-- Hex Addr	7FBB	32699
x"00",	-- Hex Addr	7FBC	32700
x"00",	-- Hex Addr	7FBD	32701
x"00",	-- Hex Addr	7FBE	32702
x"00",	-- Hex Addr	7FBF	32703
x"00",	-- Hex Addr	7FC0	32704
x"00",	-- Hex Addr	7FC1	32705
x"00",	-- Hex Addr	7FC2	32706
x"00",	-- Hex Addr	7FC3	32707
x"00",	-- Hex Addr	7FC4	32708
x"00",	-- Hex Addr	7FC5	32709
x"00",	-- Hex Addr	7FC6	32710
x"00",	-- Hex Addr	7FC7	32711
x"00",	-- Hex Addr	7FC8	32712
x"00",	-- Hex Addr	7FC9	32713
x"00",	-- Hex Addr	7FCA	32714
x"00",	-- Hex Addr	7FCB	32715
x"00",	-- Hex Addr	7FCC	32716
x"00",	-- Hex Addr	7FCD	32717
x"00",	-- Hex Addr	7FCE	32718
x"00",	-- Hex Addr	7FCF	32719
x"00",	-- Hex Addr	7FD0	32720
x"00",	-- Hex Addr	7FD1	32721
x"00",	-- Hex Addr	7FD2	32722
x"00",	-- Hex Addr	7FD3	32723
x"00",	-- Hex Addr	7FD4	32724
x"00",	-- Hex Addr	7FD5	32725
x"00",	-- Hex Addr	7FD6	32726
x"00",	-- Hex Addr	7FD7	32727
x"00",	-- Hex Addr	7FD8	32728
x"00",	-- Hex Addr	7FD9	32729
x"00",	-- Hex Addr	7FDA	32730
x"00",	-- Hex Addr	7FDB	32731
x"00",	-- Hex Addr	7FDC	32732
x"00",	-- Hex Addr	7FDD	32733
x"00",	-- Hex Addr	7FDE	32734
x"00",	-- Hex Addr	7FDF	32735
x"00",	-- Hex Addr	7FE0	32736
x"00",	-- Hex Addr	7FE1	32737
x"00",	-- Hex Addr	7FE2	32738
x"00",	-- Hex Addr	7FE3	32739
x"00",	-- Hex Addr	7FE4	32740
x"00",	-- Hex Addr	7FE5	32741
x"00",	-- Hex Addr	7FE6	32742
x"00",	-- Hex Addr	7FE7	32743
x"00",	-- Hex Addr	7FE8	32744
x"00",	-- Hex Addr	7FE9	32745
x"00",	-- Hex Addr	7FEA	32746
x"00",	-- Hex Addr	7FEB	32747
x"00",	-- Hex Addr	7FEC	32748
x"00",	-- Hex Addr	7FED	32749
x"00",	-- Hex Addr	7FEE	32750
x"00",	-- Hex Addr	7FEF	32751
x"00",	-- Hex Addr	7FF0	32752
x"00",	-- Hex Addr	7FF1	32753
x"00",	-- Hex Addr	7FF2	32754
x"00",	-- Hex Addr	7FF3	32755
x"00",	-- Hex Addr	7FF4	32756
x"00",	-- Hex Addr	7FF5	32757
x"00",	-- Hex Addr	7FF6	32758
x"00",	-- Hex Addr	7FF7	32759
x"00",	-- Hex Addr	7FF8	32760
x"00",	-- Hex Addr	7FF9	32761
x"00",	-- Hex Addr	7FFA	32762
x"00",	-- Hex Addr	7FFB	32763
x"00",	-- Hex Addr	7FFC	32764
x"00",	-- Hex Addr	7FFD	32765
x"00",	-- Hex Addr	7FFE	32766
x"00"	-- Hex Addr	7FFF	32767
);

end package;